module s1423(
  blif_clk_net,
  blif_reset_net,
  G0,
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G726,
  G729,
  G702,
  G727,
  G701BF);
input blif_clk_net;
input blif_reset_net;
input G0;
input G1;
input G2;
input G3;
input G4;
input G5;
input G6;
input G7;
input G8;
input G9;
input G10;
input G11;
input G12;
input G13;
input G14;
input G15;
input G16;
output G726;
output G729;
output G702;
output G727;
output G701BF;
reg G22;
reg G23;
reg G24;
reg G25;
reg G26;
reg G27;
reg G28;
reg G29;
reg G30;
reg G31;
reg G32;
reg G33;
reg G34;
reg G35;
reg G36;
reg G37;
reg G38;
reg G39;
reg G40;
reg G41;
reg G42;
reg G43;
reg G44;
reg G45;
reg G46;
reg G47;
reg G48;
reg G49;
reg G50;
reg G51;
reg G52;
reg G53;
reg G54;
reg G55;
reg G56;
reg G57;
reg G58;
reg G59;
reg G60;
reg G61;
reg G62;
reg G63;
reg G64;
reg G65;
reg G66;
reg G67;
reg G68;
reg G69;
reg G70;
reg G71;
reg G72;
reg G73;
reg G74;
reg G75;
reg G76;
reg G77;
reg G78;
reg G79;
reg G80;
reg G81;
reg G82;
reg G83;
reg G84;
reg G85;
reg G86;
reg G87;
reg G88;
reg G89;
reg G90;
reg G91;
reg G92;
reg G93;
reg G94;
reg G95;
wire G615;
wire G639;
wire G260;
wire G228;
wire G196;
wire G720;
wire G573;
wire G546;
wire G140;
wire G489;
wire G371;
wire G683;
wire G498;
wire G161;
wire G453;
wire G395;
wire G301;
wire G209;
wire G564;
wire G698;
wire G365;
wire G356;
wire G295;
wire G627;
wire G313;
wire G270;
wire G522;
wire G134;
wire G218;
wire G269;
wire G122;
wire G503;
wire G606;
wire G389;
wire G151;
wire G641;
wire G412;
wire G689;
wire G725;
wire G405;
wire G638;
wire G434;
wire G310;
wire II1248;
wire G238;
wire G114;
wire G302;
wire G246;
wire G175;
wire G398;
wire G172;
wire G609;
wire II1254;
wire G617;
wire G421;
wire G714;
wire G490;
wire G510;
wire G341;
wire G373;
wire G213;
wire G661;
wire G465;
wire II1242;
wire G444;
wire G716;
wire G620;
wire G354;
wire G344;
wire G300;
wire G594;
wire G722;
wire G320;
wire G566;
wire G587;
wire G488;
wire G239;
wire G419;
wire G414;
wire G312;
wire G551;
wire G227;
wire G539;
wire II1233;
wire G392;
wire G162;
wire G197;
wire G164;
wire G637;
wire G668;
wire II1267;
wire G359;
wire G364;
wire G404;
wire G141;
wire G499;
wire G123;
wire G642;
wire G343;
wire G268;
wire II1183;
wire G563;
wire G709;
wire G97;
wire G271;
wire G435;
wire G150;
wire G379;
wire G474;
wire G225;
wire G135;
wire G656;
wire G717;
wire G290;
wire G188;
wire G303;
wire G397;
wire G240;
wire G470;
wire G247;
wire G652;
wire G257;
wire G212;
wire G442;
wire G98;
wire G443;
wire G372;
wire G631;
wire G607;
wire G183;
wire G511;
wire G500;
wire G532;
wire G616;
wire G173;
wire G336;
wire G452;
wire G108;
wire G449;
wire G669;
wire G584;
wire G574;
wire G479;
wire G621;
wire G180;
wire G662;
wire G684;
wire G323;
wire G543;
wire G100;
wire G595;
wire G521;
wire G567;
wire G124;
wire G120;
wire G602;
wire G299;
wire G630;
wire G368;
wire G636;
wire G207;
wire G675;
wire G273;
wire G515;
wire G487;
wire G723;
wire G524;
wire G258;
wire G129;
wire II1;
wire G492;
wire G193;
wire G618;
wire G160;
wire G184;
wire G647;
wire G132;
wire G256;
wire G380;
wire G436;
wire G424;
wire G158;
wire G576;
wire G113;
wire G272;
wire G708;
wire G403;
wire G319;
wire G222;
wire G486;
wire II1211;
wire G558;
wire G189;
wire G592;
wire G219;
wire G441;
wire G604;
wire G338;
wire G115;
wire G480;
wire G649;
wire G417;
wire G374;
wire G243;
wire G544;
wire G157;
wire G328BF;
wire G512;
wire II1230;
wire G107;
wire G437;
wire G699;
wire G549;
wire G696;
wire G402;
wire G496;
wire G575;
wire G501;
wire G676;
wire G279;
wire G277;
wire G262;
wire G215;
wire G728;
wire G223;
wire G362;
wire G718;
wire G396;
wire G292;
wire G235;
wire G352;
wire G142;
wire G346;
wire G461;
wire G288;
wire G206;
wire G585;
wire G304;
wire G101;
wire G121;
wire G523;
wire G469;
wire G261;
wire G648;
wire G159;
wire G677;
wire G622;
wire G255;
wire G321;
wire G259;
wire G531;
wire G185;
wire G311;
wire G719;
wire G337;
wire G192;
wire G195;
wire G598;
wire G330;
wire G204;
wire G168;
wire G666;
wire G581;
wire G707;
wire G658;
wire G318;
wire G422;
wire G328;
wire G274;
wire G357;
wire G477;
wire G394;
wire G226;
wire G577;
wire G224;
wire G99;
wire G591;
wire G460;
wire G116;
wire G112;
wire G411;
wire G721;
wire G448;
wire G593;
wire G287;
wire G557;
wire G459;
wire G534;
wire G306;
wire G182;
wire G170;
wire G214;
wire G655;
wire G674;
wire G133;
wire II1257;
wire G242;
wire G440;
wire G345;
wire G550;
wire G513;
wire G401;
wire G232;
wire G686;
wire G194;
wire G605;
wire G497;
wire G667;
wire G514;
wire G278;
wire G695;
wire G701;
wire G491;
wire G305;
wire G143;
wire G429;
wire G355;
wire G472;
wire G565;
wire G106;
wire G706;
wire G178;
wire G333;
wire G381;
wire G645;
wire G167;
wire G430;
wire G234;
wire G462;
wire G291;
wire G361;
wire G590;
wire G640;
wire G138;
wire G690;
wire G438;
wire G541;
wire G623;
wire G217;
wire G200;
wire G456;
wire G353;
wire G254;
wire G191;
wire G105;
wire G144;
wire G700;
wire G670;
wire G678;
wire G329;
wire G710;
wire G147;
wire G580;
wire G493;
wire G297;
wire G117;
wire G560;
wire G506;
wire G610;
wire G447;
wire G694;
wire G600;
wire G485;
wire G176;
wire G578;
wire G210;
wire G457;
wire II1203;
wire G284;
wire G325;
wire G526;
wire G634;
wire G221;
wire G633;
wire G400;
wire G307;
wire G386;
wire G554;
wire G187;
wire G611;
wire G629;
wire G118;
wire G650;
wire G130;
wire G478;
wire G348;
wire G624;
wire G635;
wire G705;
wire G685;
wire G426;
wire G533;
wire G599;
wire G314;
wire G126;
wire G517;
wire G366;
wire G377;
wire G169;
wire G111;
wire II1227;
wire G171;
wire G263;
wire G385;
wire G233;
wire G450;
wire G324;
wire G166;
wire G507;
wire G525;
wire G446;
wire G216;
wire G471;
wire G282;
wire G286;
wire G439;
wire G369;
wire G653;
wire G145;
wire G253;
wire G596;
wire G136;
wire G494;
wire G464;
wire G332;
wire G391;
wire G190;
wire G245;
wire G155;
wire G128;
wire G409;
wire G285;
wire G308;
wire G431;
wire G420;
wire II12;
wire G603;
wire G612;
wire G688;
wire G423;
wire G559;
wire G619;
wire G316;
wire G542;
wire II1251;
wire G104;
wire G458;
wire G360;
wire G484;
wire G579;
wire G384;
wire II1245;
wire G711;
wire G205;
wire G536;
wire G375;
wire G704;
wire G673;
wire G561;
wire G376;
wire G201;
wire G264;
wire II1236;
wire G416;
wire G628;
wire G294;
wire G276;
wire G527;
wire G339;
wire II1264;
wire G509;
wire G625;
wire G547;
wire G553;
wire G127;
wire G156;
wire G657;
wire G252;
wire G332BF;
wire G110;
wire G425;
wire G475;
wire G119;
wire G131;
wire G693;
wire G516;
wire II1239;
wire G331;
wire G418;
wire G347;
wire G665;
wire G363;
wire G583;
wire G413;
wire G495;
wire G552;
wire G315;
wire G463;
wire G481;
wire G244;
wire G445;
wire G597;
wire G351;
wire G556;
wire G427;
wire G236;
wire G393;
wire G692;
wire G613;
wire G248;
wire G660;
wire G137;
wire G165;
wire G538;
wire G529;
wire G383;
wire G483;
wire G432;
wire G697;
wire G504;
wire G342;
wire G174;
wire G467;
wire G378;
wire G309;
wire G146;
wire G198;
wire G289;
wire G703;
wire G408;
wire G562;
wire G387;
wire G680;
wire G671;
wire G632;
wire G251;
wire G163;
wire G148;
wire G687;
wire G588;
wire G664;
wire G715;
wire G153;
wire G519;
wire G681;
wire G230;
wire G283;
wire G103;
wire G326;
wire G601;
wire G644;
wire G570;
wire G177;
wire G208;
wire G211;
wire G548;
wire G724;
wire G672;
wire G626;
wire G293;
wire G265;
wire G410;
wire G267;
wire G275;
wire G406;
wire G646;
wire G520;
wire G679;
wire G335;
wire G281;
wire G322;
wire G202;
wire G582;
wire G358;
wire G508;
wire G712;
wire G535;
wire II1260;
wire G370;
wire G614;
wire G149;
wire G568;
wire G468;
wire G572;
wire G713;
wire G139;
wire G109;
wire G537;
wire G237;
wire G528;
wire G555;
wire G428;
wire G473;
wire G125;
wire G691;
wire G181;
wire G659;
wire G298;
wire G454;
wire G350;
wire G476;
wire G229;
wire G296;
wire G651;
wire G199;
wire G399;
wire G482;
wire G569;
wire G589;
wire G608;
wire G179;
wire G654;
wire G502;
wire G102;
wire G317;
wire G382;
wire G388;
wire G152;
wire G643;
wire G250;
wire G241;
wire G586;
wire G334;
wire G505;
wire G407;
wire G231;
wire G280;
wire G571;
wire II1162;
wire G415;
wire G327;
wire G266;
wire G203;
wire G186;
wire G455;
wire G96;
wire G466;
wire G682;
wire G451;
wire G249;
wire G220;
wire G540;
wire G390;
wire G367;
wire G663;
wire G349;
wire G433;
wire G545;
wire G530;
wire G518;
wire G340;
wire G154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G22 <= 0;
  else
    G22 <= G332BF;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G23 <= 0;
  else
    G23 <= G328BF;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G24 <= 0;
  else
    G24 <= G109;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G25 <= 0;
  else
    G25 <= G113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G26 <= 0;
  else
    G26 <= G118;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G27 <= 0;
  else
    G27 <= G125;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G28 <= 0;
  else
    G28 <= G129;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G29 <= 0;
  else
    G29 <= G140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G30 <= 0;
  else
    G30 <= G144;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G31 <= 0;
  else
    G31 <= G149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G32 <= 0;
  else
    G32 <= G154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G33 <= 0;
  else
    G33 <= G159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G34 <= 0;
  else
    G34 <= G166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G35 <= 0;
  else
    G35 <= G175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G36 <= 0;
  else
    G36 <= G189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G37 <= 0;
  else
    G37 <= G193;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G38 <= 0;
  else
    G38 <= G198;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G39 <= 0;
  else
    G39 <= G208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G40 <= 0;
  else
    G40 <= G214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G41 <= 0;
  else
    G41 <= G218;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G42 <= 0;
  else
    G42 <= G237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G43 <= 0;
  else
    G43 <= G242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G44 <= 0;
  else
    G44 <= G247;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G45 <= 0;
  else
    G45 <= G252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G46 <= 0;
  else
    G46 <= G260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G47 <= 0;
  else
    G47 <= G303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G48 <= 0;
  else
    G48 <= G309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G49 <= 0;
  else
    G49 <= G315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G50 <= 0;
  else
    G50 <= G321;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G51 <= 0;
  else
    G51 <= G360;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G52 <= 0;
  else
    G52 <= G365;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G53 <= 0;
  else
    G53 <= G373;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G54 <= 0;
  else
    G54 <= G379;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G55 <= 0;
  else
    G55 <= G384;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G56 <= 0;
  else
    G56 <= G392;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G57 <= 0;
  else
    G57 <= G397;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G58 <= 0;
  else
    G58 <= G405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G59 <= 0;
  else
    G59 <= G408;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G60 <= 0;
  else
    G60 <= G416;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G61 <= 0;
  else
    G61 <= G424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G62 <= 0;
  else
    G62 <= G427;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G63 <= 0;
  else
    G63 <= G438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G64 <= 0;
  else
    G64 <= G441;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G65 <= 0;
  else
    G65 <= G447;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G66 <= 0;
  else
    G66 <= G451;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G67 <= 0;
  else
    G67 <= G459;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G68 <= 0;
  else
    G68 <= G464;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G69 <= 0;
  else
    G69 <= G469;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G70 <= 0;
  else
    G70 <= G477;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G71 <= 0;
  else
    G71 <= G494;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G72 <= 0;
  else
    G72 <= G498;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G73 <= 0;
  else
    G73 <= G503;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G74 <= 0;
  else
    G74 <= G526;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G75 <= 0;
  else
    G75 <= G531;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G76 <= 0;
  else
    G76 <= G536;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G77 <= 0;
  else
    G77 <= G541;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G78 <= 0;
  else
    G78 <= G548;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G79 <= 0;
  else
    G79 <= G565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G80 <= 0;
  else
    G80 <= G569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G81 <= 0;
  else
    G81 <= G573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G82 <= 0;
  else
    G82 <= G577;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G83 <= 0;
  else
    G83 <= G590;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G84 <= 0;
  else
    G84 <= G608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G85 <= 0;
  else
    G85 <= G613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G86 <= 0;
  else
    G86 <= G657;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G87 <= 0;
  else
    G87 <= G663;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G88 <= 0;
  else
    G88 <= G669;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G89 <= 0;
  else
    G89 <= G675;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G90 <= 0;
  else
    G90 <= G682;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G91 <= 0;
  else
    G91 <= G687;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G92 <= 0;
  else
    G92 <= G693;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G93 <= 0;
  else
    G93 <= G705;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G94 <= 0;
  else
    G94 <= G707;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G95 <= 0;
  else
    G95 <= G713;
assign G615 = ((~G616));
assign G639 = (G99)|(G645);
assign G260 = (G256&G258);
assign G228 = (G223&G41);
assign G196 = (G202&G37);
assign G720 = ((~II1242));
assign G573 = (G571&G572);
assign G546 = ((~G553)&(~G78));
assign G140 = (G137&G139);
assign G489 = (G508&G509);
assign G371 = ((~G372));
assign G683 = (G684&G685);
assign G498 = (G496&G497);
assign G161 = ((~G171)&(~G33));
assign G301 = ((~G50))|((~G49))|((~G48))|((~G47));
assign G209 = (G183)|(G210);
assign G453 = (G615&G445);
assign G395 = (G394&G55);
assign G564 = (G715)|(G562);
assign G698 = (G348)|(G695);
assign G365 = (G366&G364);
assign G356 = (G225)|(G355);
assign G295 = (G46)|(G105);
assign G627 = (G476)|(G645);
assign G313 = (G47)|(G311);
assign G270 = ((~G285))|((~G295));
assign G522 = (G348)|(G228);
assign G134 = (G133&G25);
assign G218 = (G219&G217);
assign G269 = ((~G284))|((~G294));
assign G122 = ((~G123))|((~G126));
assign G503 = (G501&G502);
assign G606 = (G84)|(G610);
assign G389 = ((~G395)&(~G56));
assign G151 = ((~G169)&(~G31));
assign G641 = ((~G645));
assign G412 = (G335&G57);
assign G689 = ((~G696));
assign G725 = ((~II1257));
assign G405 = (G401&G403);
assign G638 = ((~G645));
assign G434 = (G342)|(G645);
assign G310 = (G312&G313);
assign G702 = (G703&G645);
assign G238 = ((~G239)&(~G240));
assign II1248 = ((~G2));
assign G114 = ((~G115)&(~G116));
assign G302 = ((~G712));
assign G246 = ((~G259));
assign G175 = (G176&G174);
assign G398 = ((~G399)&(~G400));
assign G172 = (G171&G33);
assign G609 = ((~G610));
assign II1254 = ((~G4));
assign G617 = ((~G645));
assign G421 = ((~G431)&(~G61));
assign G714 = ((~G701));
assign G490 = (G512&G513);
assign G510 = ((~G511));
assign G341 = (G185)|(G339);
assign G373 = (G369&G371);
assign G213 = ((~G712));
assign G661 = ((~G94));
assign G465 = ((~G466)&(~G467));
assign II1242 = ((~G0));
assign G444 = ((~G615)&(~G64));
assign G716 = ((~II1230));
assign G620 = ((~G645));
assign G354 = ((~G355));
assign G344 = (G229)|(G348);
assign G300 = (G50)|(G49)|(G48)|(G47);
assign G594 = (G83)|(G593);
assign G722 = ((~II1248));
assign G320 = ((~G712));
assign G566 = ((~G610));
assign G587 = (G561)|(G78);
assign G488 = (G505&G506);
assign G239 = ((~G299)&(~G42));
assign G419 = (G358&G60);
assign G414 = (G413&G59);
assign G312 = (G48)|(G324);
assign G551 = (G550&G75);
assign G227 = (G172&G178);
assign G539 = (G551&G76);
assign II1233 = ((~G8));
assign G392 = (G388&G390);
assign G162 = (G171&G33);
assign G197 = ((~G712));
assign G164 = ((~G172))|((~G178));
assign G637 = (G722)|(G635);
assign G668 = ((~G712));
assign II1267 = ((~G95));
assign G359 = ((~G372));
assign G364 = ((~G372));
assign G404 = (G712)|(G413);
assign G141 = (G177)|(G142);
assign G499 = ((~G500));
assign G123 = ((~G135))|((~G127));
assign G642 = (G100)|(G645);
assign G343 = ((~G348));
assign G268 = ((~G288))|((~G293));
assign II1183 = ((~G11));
assign G563 = (G79)|(G610);
assign G97 = ((~G75))|((~G596));
assign G709 = (G678&G89);
assign G271 = (G275&G266);
assign G435 = (G340&G341);
assign G150 = ((~G151)&(~G152));
assign G379 = (G380&G378);
assign G474 = ((~G481)&(~G70));
assign G225 = (G204&G203);
assign G135 = (G134&G26);
assign G656 = ((~G712));
assign G717 = ((~II1233));
assign G290 = ((~G267)&(~G266));
assign G188 = ((~G712));
assign G303 = (G304&G302);
assign G397 = (G398&G396);
assign G240 = (G299&G42);
assign G470 = ((~G471)&(~G472));
assign G247 = (G248&G246);
assign G652 = (G228&G88);
assign G257 = ((~G265)&(~G46));
assign G212 = ((~G222))|((~G216));
assign G442 = ((~G443)&(~G444));
assign G98 = ((~G76))|((~G596));
assign G443 = (G615&G511);
assign G372 = (G712)|(G358);
assign G607 = (G696)|(G605);
assign G631 = (G720)|(G629);
assign G183 = (G180)|(G227);
assign G511 = ((~G63));
assign G500 = (G654)|(G712);
assign G532 = ((~G533)&(~G534));
assign G616 = ((~G482))|((~G483))|((~G484))|((~G485));
assign G452 = ((~G453)&(~G454));
assign G173 = (G172&G34);
assign G336 = ((~G355));
assign G108 = ((~G712));
assign G449 = ((~G66));
assign G669 = (G670&G668);
assign G584 = (G80)|(G75);
assign G574 = ((~G610));
assign G621 = (G614)|(G645);
assign G479 = (G434&G67);
assign G180 = ((~G92));
assign G662 = ((~G712));
assign G684 = (G645)|(G696);
assign G323 = ((~G324));
assign G543 = ((~G552)&(~G77));
assign G100 = ((~G78))|((~G596));
assign G595 = ((~G593));
assign G521 = (G487)|(G70);
assign G567 = (G80)|(G610);
assign G124 = ((~G712));
assign G120 = ((~G134)&(~G26));
assign G602 = (G85)|(G601);
assign G299 = ((~G301)&(~G328));
assign G630 = (G96)|(G645);
assign G368 = (G375&G52);
assign G636 = (G98)|(G645);
assign G207 = ((~G712));
assign G675 = (G676&G674);
assign G273 = (G278&G279);
assign G515 = ((~G72))|((~G68));
assign G487 = ((~G71)&(~G72)&(~G73));
assign G524 = (G554)|(G555);
assign G723 = ((~II1251));
assign G258 = ((~G259));
assign G129 = (G130&G128);
assign II1 = ((~G332));
assign G492 = (G71)|(G500);
assign G193 = (G194&G192);
assign G618 = (G457)|(G645);
assign G160 = ((~G161)&(~G162));
assign G184 = (G180)|(G173);
assign G647 = (G725)|(G644);
assign G256 = ((~G257)&(~G261));
assign G132 = (G136&G28);
assign G380 = ((~G381)&(~G382));
assign G436 = (G352&G353);
assign G424 = (G420&G422);
assign G158 = ((~G712));
assign G576 = (G718)|(G574);
assign G113 = (G114&G112);
assign G708 = ((~G709)&(~G710));
assign G272 = (G276&G277);
assign G403 = ((~G404));
assign G319 = (G48)|(G317);
assign G222 = (G183&G210);
assign G486 = ((~G712));
assign II1211 = ((~G701));
assign G558 = ((~G580))|((~G585));
assign G189 = (G186&G188);
assign G592 = (G594&G595);
assign G219 = ((~G220)&(~G221));
assign G441 = (G442&G440);
assign G604 = (G433&G524);
assign G338 = (G183)|(G336);
assign G115 = ((~G133)&(~G25));
assign G480 = (G479&G68);
assign G649 = (G618&G619);
assign G417 = ((~G418)&(~G419));
assign G374 = (G376&G53);
assign G243 = ((~G244)&(~G245));
assign G544 = (G552&G77);
assign G157 = (G170&G32);
assign G328BF = ((~II12));
assign G512 = (G725)|(G511);
assign G701BF = ((~II1211));
assign II1230 = ((~G7));
assign G107 = ((~G700))|((~G111));
assign G437 = ((~G712));
assign G699 = (G658)|(G712);
assign G549 = (G553&G78);
assign G696 = ((~II1203));
assign G402 = ((~G412)&(~G58));
assign G496 = (G72)|(G500);
assign G575 = (G82)|(G610);
assign G501 = (G73)|(G500);
assign G676 = (G679&G680);
assign G279 = (G268)|(G272);
assign G215 = (G222)|(G216);
assign G277 = (G267)|(G271);
assign G262 = (G299&G42);
assign G728 = ((~II1264));
assign G223 = (G222&G216);
assign G362 = ((~G523)&(~G51));
assign G718 = ((~II1236));
assign G396 = ((~G404));
assign G292 = (G43)|(G102);
assign G235 = (G649)|(G233);
assign G352 = (G346)|(G645);
assign G142 = ((~G29));
assign G346 = (G349&G350);
assign G461 = ((~G434)&(~G67));
assign G288 = ((~G44))|((~G103));
assign G206 = ((~G183))|((~G210));
assign G585 = (G81)|(G76);
assign G304 = (G306&G307);
assign G101 = (G630&G631);
assign G121 = (G134&G26);
assign G523 = (G348)|(G414);
assign G469 = (G470&G468);
assign G261 = (G265&G46);
assign G648 = (G646&G647);
assign G159 = (G160&G158);
assign G622 = (G717)|(G620);
assign G677 = ((~G678));
assign G255 = (G264&G45);
assign G321 = (G322&G320);
assign G259 = (G624&G625);
assign G531 = (G532&G530);
assign G185 = (G181&G182);
assign G311 = ((~G324));
assign G719 = ((~II1239));
assign G337 = (G224)|(G355);
assign G192 = ((~G712));
assign G195 = ((~G202)&(~G37));
assign G598 = ((~G435))|((~G83));
assign G330 = (G332&G714);
assign G204 = ((~G38));
assign G168 = (G177&G142);
assign G666 = (G87)|(G678);
assign G581 = ((~G82))|((~G77));
assign G707 = (G708&G706);
assign G658 = ((~G659));
assign G318 = (G49)|(G324);
assign G422 = ((~G423));
assign G328 = ((~G329)&(~G327));
assign G274 = (G280&G281);
assign G357 = (G184)|(G354);
assign G477 = (G473&G475);
assign G394 = (G183&G54);
assign G226 = (G136&G28);
assign G577 = (G575&G576);
assign G224 = (G203&G38);
assign G99 = ((~G77))|((~G596));
assign G591 = (G592)|(G604);
assign G460 = ((~G461)&(~G462));
assign G116 = (G133&G25);
assign G112 = ((~G712));
assign G411 = (G413&G59);
assign G721 = ((~II1245));
assign G448 = (G615)|(G65);
assign G593 = ((~G435)&(~G524));
assign G287 = ((~G43))|((~G102));
assign G557 = ((~G579))|((~G584));
assign G459 = (G460&G458);
assign G534 = (G550&G75);
assign G306 = (G47)|(G324);
assign G182 = (G35)|(G179);
assign G170 = (G169&G31);
assign G214 = (G211&G213);
assign G655 = (G91&G476);
assign G674 = ((~G712));
assign G133 = (G700&G111);
assign II1257 = ((~G5));
assign G242 = (G243&G241);
assign G440 = ((~G712));
assign G345 = (G414)|(G343);
assign G550 = (G604&G74);
assign G513 = (G722)|(G510);
assign G401 = ((~G402)&(~G406));
assign G232 = ((~G296))|((~G298))|((~G435));
assign G686 = ((~G688)&(~G660));
assign G194 = ((~G195)&(~G196));
assign G497 = (G489)|(G495);
assign G605 = ((~G610));
assign G667 = (G661)|(G665);
assign G514 = ((~G71))|((~G67));
assign G278 = (G103)|(G44);
assign G695 = ((~G696));
assign G701 = ((~G15));
assign G491 = ((~G500));
assign G305 = ((~G324));
assign G143 = ((~G712));
assign G429 = ((~G432)&(~G62));
assign G355 = (G457)|(G645);
assign G472 = (G480&G69);
assign G565 = (G563&G564);
assign G106 = ((~G107))|((~G110));
assign G706 = ((~G712));
assign G178 = ((~G34));
assign G333 = (G300)|(G714);
assign G381 = ((~G183)&(~G54));
assign G645 = ((~G90));
assign G167 = (G172)|(G178);
assign G430 = (G432&G62);
assign G234 = ((~G649))|((~G436));
assign G291 = (G42)|(G101);
assign G361 = ((~G362)&(~G363));
assign G462 = (G434&G67);
assign G590 = (G591&G588);
assign G640 = (G723)|(G638);
assign G138 = ((~G177))|((~G142));
assign G690 = (G348)|(G696);
assign G438 = (G439&G437);
assign G541 = (G542&G540);
assign G623 = ((~G645));
assign G217 = ((~G712));
assign G200 = ((~G203)&(~G38));
assign G456 = (G83)|(G524);
assign G254 = ((~G264)&(~G45));
assign G353 = (G35)|(G351);
assign G191 = ((~G36));
assign G105 = (G642&G643);
assign G144 = (G145&G143);
assign G700 = ((~G282))|((~G283));
assign G670 = (G672&G673);
assign G678 = ((~II1183));
assign G329 = (G331&G714);
assign G710 = ((~G678)&(~G94));
assign G147 = (G168&G30);
assign G580 = ((~G81))|((~G76));
assign G493 = (G488)|(G491);
assign G297 = ((~G289))|((~G290));
assign G117 = ((~G712));
assign G560 = ((~G582))|((~G587));
assign G506 = (G720)|(G504);
assign G610 = (G655)|(G712);
assign G447 = (G448&G446);
assign G485 = ((~G517))|((~G521));
assign G694 = (G697&G698);
assign G600 = ((~G601));
assign G176 = ((~G35));
assign G578 = ((~G79))|((~G74));
assign G210 = ((~G39));
assign G457 = (G455&G449&G728);
assign II1203 = ((~G10));
assign G284 = ((~G45))|((~G104));
assign G526 = (G527&G525);
assign G325 = (G50)|(G324);
assign G634 = (G721)|(G632);
assign G221 = (G223&G41);
assign G633 = (G97)|(G645);
assign G400 = (G335&G57);
assign G307 = (G719)|(G305);
assign G386 = ((~G394)&(~G55));
assign G554 = ((~G556))|((~G557))|((~G558));
assign G187 = ((~G522))|((~G191));
assign G629 = ((~G645));
assign G611 = (G85)|(G610);
assign G118 = (G119&G117);
assign G650 = (G226&G661);
assign G130 = ((~G131)&(~G132));
assign G348 = ((~G91));
assign G478 = (G481&G70);
assign G624 = (G476)|(G645);
assign G635 = ((~G645));
assign G705 = (G230&G704);
assign G685 = ((~G696));
assign G426 = ((~G712));
assign G533 = ((~G550)&(~G75));
assign G599 = ((~G598)&(~G597));
assign G126 = (G135)|(G127);
assign G314 = ((~G712));
assign G517 = ((~G487))|((~G70));
assign G366 = ((~G367)&(~G368));
assign G377 = (G183&G54&G56);
assign G169 = (G168&G30);
assign G111 = ((~G24));
assign II1227 = ((~G6));
assign G171 = (G170&G32);
assign G263 = (G262&G43);
assign G385 = ((~G386)&(~G387));
assign G233 = ((~G700))|((~G232))|((~G231));
assign G450 = ((~G712));
assign G324 = (G377)|(G348);
assign G166 = (G163&G165);
assign G507 = ((~G511));
assign G525 = ((~G589));
assign G446 = ((~G712));
assign G216 = ((~G40));
assign G471 = ((~G480)&(~G69));
assign G282 = (G105)|(G46);
assign G286 = ((~G42))|((~G101));
assign G439 = (G435)|(G63);
assign G369 = ((~G370)&(~G374));
assign G653 = (G229&G89);
assign G596 = ((~G597));
assign G145 = ((~G146)&(~G147));
assign G253 = ((~G254)&(~G255));
assign G136 = (G135&G127);
assign G494 = (G492&G493);
assign G464 = (G465&G463);
assign G332 = ((~G334))|((~G331));
assign G391 = (G712)|(G377);
assign G190 = (G522)|(G191);
assign G155 = ((~G156)&(~G157));
assign G245 = (G262&G43);
assign G128 = ((~G712));
assign G409 = ((~G410)&(~G411));
assign G285 = ((~G46))|((~G105));
assign G308 = ((~G712));
assign G420 = ((~G421)&(~G425));
assign G431 = (G358&G60);
assign II12 = ((~G328));
assign G603 = (G600)|(G84);
assign G612 = (G678)|(G609);
assign G688 = (G690&G691);
assign G423 = (G712)|(G432);
assign G559 = ((~G581))|((~G586));
assign G619 = (G715)|(G617);
assign II1251 = ((~G3));
assign G104 = (G639&G640);
assign G316 = (G318&G319);
assign G542 = ((~G543)&(~G544));
assign G458 = ((~G476));
assign G360 = (G361&G359);
assign G484 = ((~G516))|((~G520));
assign G579 = ((~G80))|((~G75));
assign G384 = (G385&G383);
assign II1245 = ((~G1));
assign G711 = ((~G712));
assign G205 = ((~G206))|((~G209));
assign G536 = (G537&G535);
assign G375 = (G523&G51);
assign G704 = ((~G712));
assign G673 = (G87)|(G671);
assign G561 = ((~G79)&(~G80)&(~G81)&(~G82));
assign G201 = (G203&G38);
assign G376 = (G375&G52);
assign II1236 = ((~G9));
assign G264 = (G263&G44);
assign G416 = (G417&G415);
assign G628 = (G718)|(G626);
assign G294 = (G45)|(G104);
assign G276 = (G102)|(G43);
assign G339 = ((~G355));
assign II1264 = ((~G16));
assign G527 = ((~G528)&(~G529));
assign G509 = (G721)|(G507);
assign G625 = (G716)|(G623);
assign G547 = ((~G589));
assign G553 = (G552&G77);
assign G127 = ((~G27));
assign G729 = ((~II1267));
assign G156 = ((~G170)&(~G32));
assign G657 = (G659&G656);
assign G252 = (G253&G251);
assign G110 = (G700)|(G111);
assign G332BF = ((~II1));
assign G425 = (G431&G61);
assign G475 = ((~G476));
assign G119 = ((~G120)&(~G121));
assign G131 = ((~G136)&(~G28));
assign G693 = (G692)|(G699);
assign G516 = ((~G73))|((~G69));
assign II1239 = ((~G12));
assign G331 = ((~G333))|((~G22));
assign G418 = ((~G358)&(~G60));
assign G347 = ((~G348));
assign G665 = ((~G678));
assign G363 = (G523&G51);
assign G583 = (G79)|(G74);
assign G495 = ((~G500));
assign G413 = (G335&G58);
assign G552 = (G551&G76);
assign G315 = (G316&G314);
assign G463 = ((~G476));
assign G481 = (G480&G69);
assign G244 = ((~G262)&(~G43));
assign G597 = ((~G602))|((~G603));
assign G445 = ((~G65));
assign G351 = ((~G645));
assign G556 = ((~G578))|((~G583));
assign G427 = (G428&G426);
assign G236 = ((~G259));
assign G692 = ((~G694)&(~G660));
assign G393 = (G395&G56);
assign G613 = (G611&G612);
assign G248 = ((~G249)&(~G250));
assign G660 = ((~G658)&(~G86));
assign G137 = ((~G138))|((~G141));
assign G165 = ((~G712));
assign G538 = ((~G551)&(~G76));
assign G383 = ((~G391));
assign G529 = (G604&G74);
assign G483 = ((~G515))|((~G519));
assign G432 = (G358&G61);
assign G697 = (G180)|(G696);
assign G504 = ((~G511));
assign G174 = ((~G712));
assign G342 = (G344&G345);
assign G467 = (G479&G68);
assign G146 = ((~G168)&(~G30));
assign G378 = ((~G391));
assign G309 = (G310&G308);
assign G198 = (G199&G197);
assign G289 = ((~G270)&(~G269)&(~G268));
assign G703 = ((~G650)&(~G651)&(~G652)&(~G653));
assign G408 = (G409&G407);
assign G562 = ((~G610));
assign G387 = (G394&G55);
assign G680 = (G88)|(G677);
assign G671 = ((~G678));
assign G632 = ((~G645));
assign G251 = ((~G259));
assign G163 = ((~G164))|((~G167));
assign G148 = ((~G712));
assign G588 = ((~G589));
assign G687 = (G686)|(G699);
assign G715 = ((~II1227));
assign G664 = (G666&G667);
assign G153 = ((~G712));
assign G519 = (G72)|(G68);
assign G681 = ((~G683)&(~G660));
assign G230 = ((~G234))|((~G235));
assign G283 = (G270)|(G274);
assign G727 = (G476&G645);
assign G103 = (G636&G637);
assign G601 = (G621&G622);
assign G326 = (G49)|(G323);
assign G644 = ((~G645));
assign G570 = ((~G610));
assign G177 = (G180)|(G226);
assign G208 = (G205&G207);
assign G724 = ((~II1254));
assign G548 = (G545&G547);
assign G211 = ((~G212))|((~G215));
assign G672 = (G88)|(G678);
assign G626 = ((~G645));
assign G293 = (G44)|(G103);
assign G265 = (G264&G45);
assign G410 = ((~G413)&(~G59));
assign G267 = ((~G287))|((~G292));
assign G275 = (G101)|(G42);
assign G406 = (G412&G58);
assign G646 = (G456)|(G645);
assign G520 = (G73)|(G69);
assign G679 = (G89)|(G678);
assign G335 = (G337&G338);
assign G281 = (G269)|(G273);
assign G322 = (G325&G326);
assign G202 = (G522&G191);
assign G582 = ((~G561))|((~G78));
assign G358 = (G523&G53);
assign G508 = (G724)|(G511);
assign G712 = ((~G14));
assign G535 = ((~G589));
assign II1260 = ((~G93));
assign G370 = ((~G376)&(~G53));
assign G614 = ((~G64));
assign G149 = (G150&G148);
assign G568 = (G716)|(G566);
assign G468 = ((~G476));
assign G572 = (G717)|(G570);
assign G713 = (G599&G711);
assign G139 = ((~G712));
assign G109 = (G106&G108);
assign G537 = ((~G538)&(~G539));
assign G237 = (G238&G236);
assign G528 = ((~G604)&(~G74));
assign G555 = ((~G559))|((~G560));
assign G428 = ((~G429)&(~G430));
assign G473 = ((~G474)&(~G478));
assign G125 = (G122&G124);
assign G691 = (G645)|(G689);
assign G659 = ((~II1162));
assign G181 = (G178)|(G180);
assign G298 = ((~G297))|((~G700));
assign G454 = ((~G615)&(~G66));
assign G476 = ((~G486))|((~G616));
assign G350 = (G59)|(G347);
assign G229 = (G432&G62);
assign G296 = ((~G297));
assign G199 = ((~G200)&(~G201));
assign G651 = (G227&G87);
assign G399 = ((~G335)&(~G57));
assign G482 = ((~G514))|((~G518));
assign G569 = (G567&G568);
assign G589 = (G627&G628);
assign G608 = (G606&G607);
assign G179 = ((~G180));
assign G654 = (G90&G476);
assign G102 = (G633&G634);
assign G502 = (G490)|(G499);
assign G317 = ((~G324));
assign G152 = (G169&G31);
assign G382 = (G183&G54);
assign G388 = ((~G389)&(~G393));
assign G643 = (G724)|(G641);
assign G250 = (G263&G44);
assign G241 = ((~G259));
assign G586 = (G82)|(G77);
assign G334 = (G301)|(G714);
assign G407 = ((~G712));
assign G505 = (G723)|(G511);
assign G231 = ((~G435))|((~G648));
assign II1162 = ((~G13));
assign G280 = (G104)|(G45);
assign G571 = (G81)|(G610);
assign G415 = ((~G423));
assign G327 = ((~G330)&(~G23));
assign G266 = ((~G286))|((~G291));
assign G455 = ((~G456));
assign G186 = ((~G187))|((~G190));
assign G203 = (G202&G37);
assign G96 = ((~G74))|((~G596));
assign G466 = ((~G479)&(~G68));
assign G682 = (G681)|(G699);
assign G451 = (G452&G450);
assign G249 = ((~G263)&(~G44));
assign G220 = ((~G223)&(~G41));
assign G540 = ((~G589));
assign G390 = ((~G391));
assign G367 = ((~G375)&(~G52));
assign G663 = (G664&G662);
assign G349 = (G62)|(G348);
assign G433 = (G356&G357);
assign G545 = ((~G546)&(~G549));
assign G530 = ((~G589));
assign G518 = (G71)|(G67);
assign G154 = (G155&G153);
assign G340 = (G38)|(G355);
assign G726 = ((~II1260));
endmodule
