module s386(
  blif_clk_net,
  blif_reset_net,
  v6,
  v5,
  v4,
  v3,
  v2,
  v1,
  v0,
  v13_D_12,
  v13_D_11,
  v13_D_10,
  v13_D_9,
  v13_D_8,
  v13_D_7,
  v13_D_6);
input blif_clk_net;
input blif_reset_net;
input v6;
input v5;
input v4;
input v3;
input v2;
input v1;
input v0;
output v13_D_12;
output v13_D_11;
output v13_D_10;
output v13_D_9;
output v13_D_8;
output v13_D_7;
output v13_D_6;
reg v12;
reg v11;
reg v10;
reg v9;
reg v8;
reg v7;
wire B30B;
wire IIII102;
wire II158;
wire IIII108;
wire Lv13_D_3;
wire IIII71;
wire Lv13_D_5;
wire IIII25;
wire II195;
wire II207;
wire B31B;
wire B42B;
wire IIII27;
wire II175;
wire II222;
wire IIII100;
wire B44B;
wire IIII39;
wire IIII28;
wire Lv13_D_9;
wire II64;
wire IIII77;
wire II124;
wire B45B;
wire IIII93;
wire Lv13_D_11;
wire IIII57;
wire IIII73;
wire IIII106;
wire IIII18;
wire IIII62;
wire Lv13_D_7;
wire B34Bbar;
wire IIII31;
wire II167;
wire B16B;
wire B29B;
wire IIII69;
wire IIII113;
wire IIII43;
wire v13_D_4;
wire II231;
wire B40B;
wire B26B;
wire IIII63;
wire II225;
wire IIII41;
wire v13_D_2;
wire v13_D_1;
wire IIII66;
wire B35Bbar;
wire IIII48;
wire v3bar;
wire Lv13_D_1;
wire IIII84;
wire II98;
wire IIII47;
wire B35B;
wire II148;
wire IIII22;
wire B38B;
wire B32B;
wire IIII74;
wire B19B;
wire B28B;
wire II171;
wire B23B;
wire Lv13_D_10;
wire II204;
wire v6bar;
wire IIII51;
wire IIII90;
wire II213;
wire B25B;
wire IIII53;
wire II89;
wire IIII96;
wire II210;
wire v7bar;
wire B36B;
wire v13_D_0;
wire B18B;
wire v12bar;
wire II234;
wire v0bar;
wire Lv13_D_2;
wire IIII98;
wire IIII35;
wire II104;
wire IIII87;
wire IIII54;
wire B15B;
wire v11bar;
wire IIII76;
wire B27B;
wire II201;
wire II97;
wire II198;
wire II65;
wire B43B;
wire IIII105;
wire II216;
wire IIII59;
wire B20B;
wire B39B;
wire B37B;
wire II228;
wire B14B;
wire v4bar;
wire IIII111;
wire B14Bbar;
wire Lv13_D_6;
wire IIII24;
wire B17B;
wire IIII30;
wire IIII17;
wire IIII36;
wire Lv13_D_4;
wire IIII103;
wire B33B;
wire B21B;
wire B24B;
wire IIII44;
wire v8bar;
wire IIII85;
wire IIII109;
wire v1bar;
wire v13_D_3;
wire B34B;
wire B22B;
wire IIII94;
wire IIII65;
wire IIII21;
wire II186;
wire Lv13_D_0;
wire Lv13_D_12;
wire II192;
wire IIII60;
wire IIII91;
wire Lv13_D_8;
wire IIII50;
wire IIII114;
wire II219;
wire IIII40;
wire II164;
wire IIII56;
wire v10bar;
wire IIII79;
wire B41B;
wire v9bar;
wire v13_D_5;
wire v5bar;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v12 <= 0;
  else
    v12 <= v13_D_5;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v11 <= 0;
  else
    v11 <= v13_D_4;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v10 <= 0;
  else
    v10 <= v13_D_3;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v9 <= 0;
  else
    v9 <= v13_D_2;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v8 <= 0;
  else
    v8 <= v13_D_1;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v7 <= 0;
  else
    v7 <= v13_D_0;
assign B30B = (IIII71)|(v7);
assign IIII102 = (v8bar&v11bar&v12);
assign II158 = (B39B&v7bar&v9bar);
assign IIII108 = (v7&v11);
assign v13_D_7 = ((~II213));
assign Lv13_D_3 = (IIII35)|(IIII36);
assign IIII71 = (v4bar&v11bar&B34Bbar);
assign Lv13_D_5 = (v9bar&v10bar&II167);
assign IIII25 = (v0bar&B22B);
assign II195 = (B20B&v0&v1bar);
assign II207 = ((~Lv13_D_9));
assign v13_D_12 = ((~II198));
assign B31B = (IIII43)|(IIII44);
assign B42B = (IIII111)|(v12bar);
assign IIII27 = (B44B&v10bar);
assign II175 = (v0&v7bar&v8bar);
assign II222 = ((~Lv13_D_4));
assign IIII100 = (v2&v8bar);
assign B44B = (IIII59)|(IIII60);
assign IIII39 = (v5&v7&v8bar&v11);
assign IIII28 = (v10&v11bar&v12bar&II175);
assign Lv13_D_9 = (v11bar&v12bar&II158);
assign II64 = (v0bar&v5&v7bar&v8bar);
assign IIII77 = (v0&v8bar&v10);
assign II124 = (B40B&v1&v7bar&v8bar);
assign B45B = (IIII27)|(IIII28);
assign IIII93 = (v9bar&v10bar);
assign Lv13_D_11 = (IIII17)|(IIII18);
assign IIII57 = (B32B&v7bar);
assign IIII73 = (v4bar&v11bar&B34Bbar);
assign IIII106 = (v5bar&v7bar&v11&v12);
assign IIII18 = (v0bar&v10bar&B41B);
assign IIII62 = (B23B&v7bar&v8bar);
assign Lv13_D_7 = (v9bar&v10bar&v12bar&II148);
assign B34Bbar = ((~B34B));
assign IIII31 = (B36B&v11bar&v12bar);
assign II167 = (B33B&v0&v1bar);
assign B16B = (B35Bbar)|(IIII69);
assign B29B = (IIII105)|(IIII106);
assign IIII69 = (v7&v11bar);
assign IIII113 = (v7bar&v8bar);
assign IIII43 = (B30B&v12bar);
assign v13_D_4 = ((~II222));
assign II231 = ((~Lv13_D_1));
assign B40B = (IIII98)|(v10bar);
assign B26B = (v0bar)|(IIII96);
assign IIII63 = (v9bar&v10bar&v12bar);
assign II225 = ((~Lv13_D_3));
assign IIII41 = (v4&v11bar&B17B);
assign v13_D_1 = ((~II231));
assign v13_D_2 = ((~II228));
assign v13_D_11 = ((~II201));
assign IIII66 = (v4&v7);
assign B35Bbar = ((~B35B));
assign IIII48 = (B14B&v11);
assign v3bar = ((~v3));
assign Lv13_D_1 = (v9bar&v10bar&II195);
assign IIII84 = (v8bar&v11&v12);
assign II98 = (v9bar&v10&v11bar&v12bar);
assign IIII47 = (v4bar&v11bar&B34Bbar);
assign B35B = (v2)|(v7);
assign II148 = (B38B&v0&v1bar);
assign IIII22 = (v7bar&B18B);
assign B38B = (IIII73)|(IIII74);
assign B32B = (IIII84)|(IIII85);
assign IIII74 = (v7&v8bar&v11);
assign B19B = (IIII39)|(IIII40)|(IIII41);
assign B28B = (IIII53)|(IIII54);
assign II171 = (v5&v7bar&v8bar);
assign B23B = (IIII90)|(IIII91);
assign Lv13_D_10 = (v9&v11bar&v12bar&II124);
assign II204 = ((~Lv13_D_10));
assign v6bar = ((~v6));
assign IIII51 = (v9bar&v10bar&v12bar);
assign IIII90 = (v9bar&v10bar);
assign II213 = ((~Lv13_D_7));
assign B25B = (v10bar)|(IIII79);
assign IIII53 = (B27B&v1);
assign II89 = (v5bar&v7bar&v8bar);
assign IIII96 = (v1&v9bar);
assign II210 = ((~Lv13_D_8));
assign v13_D_6 = ((~II216));
assign v7bar = ((~v7));
assign B36B = (IIII65)|(IIII66);
assign v13_D_0 = ((~II234));
assign B18B = (IIII102)|(IIII103);
assign v12bar = ((~v12));
assign v0bar = ((~v0));
assign II234 = ((~Lv13_D_0));
assign Lv13_D_2 = (IIII24)|(IIII25);
assign IIII98 = (v0&v5);
assign IIII35 = (B28B&v12bar);
assign II104 = (v2&v3&v8);
assign IIII87 = (v5bar&v9&v11bar&v12bar);
assign IIII54 = (v0bar&v9bar&v10bar);
assign B15B = (IIII47)|(IIII48);
assign v11bar = ((~v11));
assign IIII76 = (v1bar&v4&v10bar&B34Bbar);
assign v13_D_8 = ((~II210));
assign II201 = ((~Lv13_D_11));
assign II97 = (v0&v6bar&v7bar&v8bar);
assign B27B = (IIII93)|(IIII94);
assign II198 = ((~Lv13_D_12));
assign II65 = (v9&v10&v11bar&v12bar);
assign B43B = (IIII108)|(IIII109);
assign IIII105 = (v2&v11bar&v12bar);
assign II216 = ((~Lv13_D_6));
assign IIII59 = (B43B&v8&v12bar);
assign B20B = (IIII21)|(IIII22);
assign B39B = (IIII76)|(IIII77);
assign B37B = (IIII30)|(IIII31);
assign II228 = ((~Lv13_D_2));
assign B14B = (v7bar)|(v8bar);
assign v4bar = ((~v4));
assign IIII111 = (v7bar&v8bar);
assign IIII24 = (B24B&v1);
assign B14Bbar = ((~B14B));
assign Lv13_D_6 = (v9bar&v10bar&II192);
assign B17B = (v7)|(IIII100);
assign IIII17 = (B45B&v9bar);
assign IIII30 = (v11&v12&II171);
assign IIII36 = (v7bar&v8bar&B25B&B26B);
assign Lv13_D_4 = (v9bar&v10bar&II186);
assign v13_D_10 = ((~II204));
assign IIII103 = (v8&v11&v12bar);
assign B33B = (IIII56)|(IIII57);
assign B21B = (v10bar)|(IIII87);
assign B24B = (IIII62)|(IIII63);
assign v8bar = ((~v8));
assign IIII44 = (v8bar&B29B);
assign IIII85 = (v11bar&v12bar&II104);
assign IIII109 = (v3bar&v4bar&v11bar);
assign v1bar = ((~v1));
assign v13_D_3 = ((~II225));
assign B34B = (v8bar)|(v3);
assign B22B = (IIII50)|(IIII51);
assign IIII94 = (v10&v11bar&II89);
assign IIII65 = (B35B&B34B);
assign IIII21 = (B19B&v12bar);
assign II186 = (B31B&v0&v1bar);
assign Lv13_D_0 = (v9bar&v10bar&v12bar&II164);
assign Lv13_D_12 = (II64&II65);
assign II192 = (B37B&v0&v1bar);
assign IIII60 = (v1&B42B);
assign IIII91 = (v0&v11bar&v12bar);
assign Lv13_D_8 = (II97&II98);
assign IIII50 = (B21B&v7bar&v8bar);
assign IIII114 = (v9bar&v12bar);
assign v13_D_9 = ((~II207));
assign II219 = ((~Lv13_D_5));
assign II164 = (B15B&v0&v1bar);
assign IIII40 = (v3&v8&B16B);
assign IIII56 = (v11&v12bar&B14Bbar);
assign v10bar = ((~v10));
assign IIII79 = (v11bar&v12bar);
assign B41B = (IIII113)|(IIII114);
assign v13_D_5 = ((~II219));
assign v9bar = ((~v9));
assign v5bar = ((~v5));
endmodule
