module s510(
  blif_clk_net,
  blif_reset_net,
  john,
  cnt13,
  cnt21,
  cnt284,
  pcnt6,
  cnt261,
  cnt44,
  pcnt12,
  pcnt17,
  cnt591,
  cnt45,
  cnt567,
  pcnt27,
  cnt283,
  cnt272,
  cnt10,
  cnt511,
  pcnt241,
  cnt509,
  csm,
  pclr,
  pc,
  cclr,
  vsync,
  cblank,
  csync);
input blif_clk_net;
input blif_reset_net;
input john;
input cnt13;
input cnt21;
input cnt284;
input pcnt6;
input cnt261;
input cnt44;
input pcnt12;
input pcnt17;
input cnt591;
input cnt45;
input cnt567;
input pcnt27;
input cnt283;
input cnt272;
input cnt10;
input cnt511;
input pcnt241;
input cnt509;
output csm;
output pclr;
output pc;
output cclr;
output vsync;
output cblank;
output csync;
reg st_5;
reg st_4;
reg st_3;
reg st_2;
reg st_1;
reg st_0;
wire II798;
wire II739;
wire II539;
wire II909_1;
wire II1102_1;
wire II855;
wire II924_1;
wire II1116_2;
wire II1062_1;
wire II946_2;
wire II663;
wire II872;
wire II207;
wire II209;
wire II574;
wire II494;
wire II978_1;
wire II535;
wire II547;
wire II595;
wire II326;
wire II587;
wire II531;
wire II731;
wire II810;
wire II1077_1;
wire II95;
wire II958_2;
wire II130;
wire II270;
wire II921_1;
wire II495;
wire II591;
wire II7;
wire II823;
wire II943_1;
wire II936_1;
wire II1110_1;
wire II779;
wire II877;
wire II486;
wire II6;
wire II874;
wire II1074_1;
wire II615;
wire II506;
wire II1089_1;
wire II936_2;
wire II59;
wire II131;
wire II70;
wire II889;
wire II266;
wire II232;
wire II1106_1;
wire II1123_1;
wire II474;
wire II60;
wire II4;
wire II903_2;
wire II861;
wire II1085_2;
wire II782;
wire II217;
wire II863;
wire II478;
wire II954_2;
wire II278;
wire II1055_2;
wire II710;
wire II928_1;
wire II466;
wire II68;
wire II962_2;
wire II787;
wire II917_2;
wire II1085_1;
wire II837;
wire II1099_1;
wire II487;
wire II841;
wire II982_1;
wire II1044_1;
wire II627;
wire II774;
wire II583;
wire II638;
wire II462;
wire II642;
wire II511;
wire II940_1;
wire II78;
wire II946_1;
wire II230;
wire II259;
wire II204;
wire II950_1;
wire II671;
wire II58;
wire II213;
wire II67;
wire II988_1;
wire II607;
wire II924_2;
wire II543;
wire II1071_1;
wire II618;
wire II814;
wire II1102_2;
wire II555;
wire II498;
wire II347;
wire II887;
wire II1095_2;
wire II903_1;
wire II234;
wire II658;
wire II1065_1;
wire II958_1;
wire II598;
wire II867;
wire II490;
wire II747;
wire II104;
wire II698;
wire II551;
wire II714;
wire II667;
wire II458;
wire II1116_1;
wire II371;
wire II675;
wire II834;
wire II216;
wire II298;
wire II578;
wire II56;
wire II69;
wire II390;
wire II603;
wire II566;
wire II917_1;
wire II821;
wire II546;
wire II881;
wire II73;
wire II962_1;
wire II5;
wire II666;
wire II827;
wire II274;
wire II594;
wire II2;
wire II795;
wire II282;
wire II778;
wire II1081_2;
wire II1092_1;
wire II985_1;
wire II1120_1;
wire II590;
wire II475;
wire II570;
wire II799;
wire II1038_1;
wire II884;
wire II57;
wire II1055_1;
wire II1113_1;
wire II563;
wire II899;
wire II205;
wire II1106_2;
wire II933_1;
wire II1059_1;
wire II838;
wire II954_1;
wire II61;
wire II914_1;
wire II455;
wire II559;
wire II467;
wire II1068_1;
wire II1081_1;
wire II1095_1;
wire II900_1;
wire II554;
wire II463;
wire II742;
wire II975_1;
wire II346;
wire II950_2;
wire II895;
wire II567;
wire II967_1;
wire II530;
wire II831;
wire II970_1;
wire II482;
wire II3;
wire II483;
wire II694;
wire II870;
wire II606;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    st_5 <= 0;
  else
    st_5 <= II2;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    st_4 <= 0;
  else
    st_4 <= II3;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    st_3 <= 0;
  else
    st_3 <= II4;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    st_2 <= 0;
  else
    st_2 <= II5;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    st_1 <= 0;
  else
    st_1 <= II6;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    st_0 <= 0;
  else
    st_0 <= II7;
assign II798 = ((~II799));
assign II739 = ((~st_5)&(~st_1));
assign II909_1 = (II466)|(II627);
assign II539 = ((~II546)&(~II60));
assign II1102_1 = (st_5&II455);
assign II855 = ((~II615)&(~st_3));
assign vsync = ((~II914_1))|((~II855))|((~II867));
assign II924_1 = (st_0)|(II731);
assign II1116_2 = (II61&II230);
assign II1062_1 = (II535&II598);
assign II663 = ((~st_1)&(~II58));
assign II946_2 = (john&st_4);
assign II872 = ((~II1095_1))|((~II1095_2))|((~II774));
assign II207 = ((~II595)&(~II943_1));
assign II574 = ((~st_3))|((~II57));
assign II209 = ((~II946_1)&(~II946_2));
assign II494 = ((~II57))|((~II547));
assign II978_1 = (II483)|(II747);
assign II535 = ((~II590)&(~st_0));
assign II547 = ((~II61)&(~st_2));
assign II595 = ((~st_0)&(~st_2));
assign II326 = ((~II982_1))|((~II61));
assign II587 = ((~st_1)&(~st_2));
assign II531 = ((~II574)&(~II59));
assign II731 = ((~II583)&(~II607));
assign II810 = ((~pcnt6))|((~cnt284))|((~II455));
assign II1077_1 = (II104&II539);
assign II95 = ((~II587)&(~II591));
assign II958_2 = (cnt284)|(II642);
assign cclr = ((~II486))|((~II877))|((~II546))|((~II390));
assign II270 = ((~st_3))|((~II615));
assign II921_1 = (II494)|(II570);
assign II130 = ((~II131));
assign II495 = ((~II494));
assign II7 = ((~II778))|((~II782))|((~II887));
assign II591 = ((~II590));
assign II823 = ((~II259)&(~II1059_1));
assign pclr = ((~II917_1))|((~II917_2));
assign II943_1 = (II578&st_3);
assign II936_1 = (cnt591&II59);
assign II1110_1 = (II61)|(II530);
assign II779 = ((~II95)&(~st_4)&(~II638));
assign II877 = ((~II1102_1)&(~II1102_2)&(~II551));
assign II486 = ((~II487));
assign csm = ((~II555)&(~II798));
assign II6 = ((~II909_1))|((~II899))|((~II895));
assign II874 = ((~II1099_1))|((~II863))|((~II831));
assign II1074_1 = (II475)|(II546);
assign II615 = ((~II475)&(~st_2));
assign II506 = ((~II535))|((~II58));
assign II1089_1 = (II59&II555);
assign II936_2 = (cnt272&st_2);
assign cblank = ((~II928_1))|((~II841));
assign II59 = ((~st_2));
assign II131 = ((~II936_1)&(~II936_2));
assign II70 = ((~pcnt17));
assign II889 = ((~II1116_1)&(~II1116_2)&(~II870));
assign II266 = ((~II970_1))|((~st_1));
assign II232 = ((~II962_1))|((~II962_2))|((~II810));
assign II1106_1 = (II60&II551);
assign II1123_1 = (II551&II663);
assign II60 = ((~st_1));
assign II474 = ((~II56))|((~II57));
assign II903_2 = (II58)|(II478);
assign II4 = ((~II278))|((~II274))|((~II270))|((~II266));
assign II861 = ((~II1081_1)&(~II1081_2));
assign II1085_2 = (II61&II216);
assign II782 = ((~II67))|((~II559))|((~II675));
assign II217 = ((~II954_1)&(~II954_2));
assign II863 = ((~II1085_1)&(~II1085_2));
assign II478 = ((~II547))|((~II739));
assign II954_2 = (cnt45&II587&II104);
assign II278 = ((~II975_1))|((~II60));
assign II710 = ((~II467))|((~cnt10));
assign II1055_2 = (II58&II204);
assign II928_1 = (st_0)|(II530);
assign II466 = ((~st_3))|((~II535));
assign II68 = ((~cnt44));
assign II962_2 = (II466)|(II78);
assign II787 = ((~II554)&(~st_5)&(~II574));
assign II917_2 = (II482)|(II590);
assign II837 = ((~II487)&(~II1071_1));
assign II1085_1 = (II787&II130);
assign II1099_1 = (II506)|(II209);
assign II487 = ((~st_4)&(~II498));
assign II841 = ((~II799)&(~II1077_1));
assign II982_1 = (II559)|(II487);
assign II1044_1 = (II70&cnt284);
assign II627 = ((~pcnt241)&(~II78));
assign II583 = ((~II511)&(~II60));
assign II774 = ((~st_5))|((~II547))|((~II458));
assign II638 = ((~II511))|((~st_0));
assign II462 = ((~II463));
assign II511 = ((~st_3)&(~st_5));
assign II642 = ((~II739))|((~st_2));
assign II940_1 = (II495&II60);
assign II78 = ((~cnt511));
assign II946_1 = (cnt10&st_5);
assign II230 = ((~II958_1))|((~II958_2));
assign II259 = ((~st_0)&(~II967_1));
assign II204 = ((~II205));
assign II950_1 = (II455&cnt45);
assign II671 = ((~II458)&(~II59));
assign II58 = ((~st_3));
assign II213 = ((~II950_1)&(~II950_2));
assign II67 = ((~cnt261));
assign II924_2 = (II474)|(II666);
assign II988_1 = (II694&II698);
assign II607 = ((~II606));
assign II543 = ((~II742)&(~II590));
assign II1071_1 = (II551&II671);
assign II618 = ((~II69))|((~cnt44));
assign II814 = ((~II58))|((~cnt21))|((~II595));
assign II1102_2 = (II56&II675);
assign II555 = ((~st_0)&(~st_1));
assign II498 = ((~II511))|((~II587));
assign II347 = ((~II346));
assign II887 = ((~II874)&(~II1113_1));
assign II1095_2 = (II475)|(II578);
assign II903_1 = (II606)|(II742);
assign II234 = ((~II213))|((~II814))|((~II710))|((~II714));
assign II658 = ((~st_2))|((~II58));
assign II1065_1 = (II475&II232);
assign II958_1 = (II57)|(II59);
assign II598 = ((~cnt13))|((~II56));
assign II867 = ((~II834)&(~II1089_1));
assign II490 = ((~cnt284))|((~pcnt17));
assign II747 = ((~II638)&(~II1044_1));
assign II104 = ((~II933_1))|((~II56));
assign II551 = ((~II61)&(~II57));
assign II698 = ((~II563))|((~II59));
assign II714 = ((~II1038_1))|((~II567));
assign II667 = ((~II666));
assign II458 = ((~st_3))|((~st_1));
assign II1116_1 = (II95&II603);
assign II371 = ((~II68)&(~II988_1));
assign II675 = ((~II61)&(~st_1));
assign II834 = ((~II1068_1))|((~II642));
assign II298 = ((~II539))|((~II574));
assign II216 = ((~II217));
assign II578 = ((~II61))|((~st_1));
assign II56 = ((~st_5));
assign II69 = ((~pcnt12));
assign II390 = ((~st_0))|((~II583));
assign pc = ((~II921_1))|((~II837));
assign II603 = ((~II61)&(~II56));
assign II566 = ((~II663))|((~st_2));
assign II821 = ((~II1055_1)&(~II1055_2));
assign II917_1 = (II458)|(II494)|(st_5);
assign II881 = ((~II1106_1)&(~II1106_2)&(~II838));
assign II546 = ((~II547));
assign II73 = ((~cnt567));
assign II962_1 = (II462)|(II73);
assign II666 = ((~II61))|((~st_3));
assign II5 = ((~II282))|((~II889))|((~II827))|((~II298));
assign II827 = ((~II531)&(~II1062_1));
assign II274 = ((~II56))|((~II667));
assign II594 = ((~II595));
assign csync = ((~II924_1))|((~II924_2))|((~II881));
assign II2 = ((~II900_1))|((~II821));
assign II282 = ((~II978_1))|((~st_1));
assign II795 = ((~st_3)&(~st_2)&(~II578));
assign II778 = ((~II779));
assign II1081_2 = (st_2&II483);
assign II985_1 = (pcnt27)|(II73);
assign II1092_1 = (st_4)|(II478);
assign II590 = ((~st_1))|((~st_2));
assign II475 = ((~II474));
assign II1120_1 = (II795&II618);
assign II570 = ((~II458))|((~II56));
assign II799 = ((~II56)&(~II58)&(~II59));
assign II1038_1 = (cnt21)|(st_0);
assign II884 = ((~II1110_1))|((~II861))|((~II326));
assign II57 = ((~st_4));
assign II1055_1 = (II570&st_0&st_2);
assign II563 = ((~II578)&(~II56));
assign II1113_1 = (st_4&II234);
assign II899 = ((~II872)&(~II347)&(~II1123_1));
assign II205 = ((~II563)&(~II940_1));
assign II1106_2 = (II57&II543);
assign II933_1 = (II57)|(II58);
assign II1059_1 = (st_5&II671);
assign II838 = ((~II1074_1))|((~II530));
assign II61 = ((~st_0));
assign II954_1 = (st_5&cnt509&II567);
assign II914_1 = (II60)|(II61);
assign II455 = ((~II554)&(~II658));
assign II559 = ((~II658)&(~II56));
assign II467 = ((~II466));
assign II1081_1 = (II543&II490&II58);
assign II1068_1 = (st_4)|(II590);
assign II1095_1 = (cnt13)|(II506);
assign II900_1 = (II56)|(II207);
assign II554 = ((~II555));
assign II463 = ((~II458)&(~II594));
assign II742 = ((~II56))|((~st_0));
assign II975_1 = (II531)|(II483);
assign II346 = ((~II985_1))|((~II463));
assign II950_2 = (II463&cnt283);
assign II895 = ((~II884)&(~II1120_1));
assign II567 = ((~II566));
assign II967_1 = (II498&II57);
assign II530 = ((~II531));
assign II831 = ((~II371)&(~II1065_1));
assign II970_1 = (II495)|(II603);
assign II482 = ((~II58))|((~II551));
assign II3 = ((~II903_1))|((~II903_2))|((~II823));
assign II483 = ((~II482));
assign II694 = ((~II795))|((~II57));
assign II870 = ((~II1092_1))|((~II566));
assign II606 = ((~II95))|((~II57));
endmodule
