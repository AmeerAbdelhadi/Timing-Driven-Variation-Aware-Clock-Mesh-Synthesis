module s1196(
  blif_clk_net,
  blif_reset_net,
  G0,
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G546,
  G539,
  G550,
  G551,
  G552,
  G547,
  G548,
  G549,
  G530,
  G45,
  G542,
  G532,
  G535,
  G537);
input blif_clk_net;
input blif_reset_net;
input G0;
input G1;
input G2;
input G3;
input G4;
input G5;
input G6;
input G7;
input G8;
input G9;
input G10;
input G11;
input G12;
input G13;
output G546;
output G539;
output G550;
output G551;
output G552;
output G547;
output G548;
output G549;
output G530;
output G45;
output G542;
output G532;
output G535;
output G537;
reg G29;
reg G30;
reg G31;
reg G32;
reg G33;
reg G34;
reg G35;
reg G36;
reg G37;
reg G38;
reg G39;
reg G40;
reg G41;
reg G42;
reg G43;
reg G44;
reg G45;
reg G46;
wire G260;
wire G228;
wire G196;
wire G61;
wire G140;
wire G371;
wire G489;
wire G498;
wire G161;
wire G395;
wire G209;
wire G301;
wire G453;
wire G365;
wire G356;
wire G295;
wire G313;
wire G270;
wire G522;
wire G218;
wire G134;
wire G269;
wire G83;
wire G80;
wire G122;
wire G503;
wire G389;
wire G151;
wire G412;
wire G405;
wire G81;
wire G58;
wire G434;
wire G310;
wire G238;
wire G114;
wire II218;
wire G302;
wire G246;
wire G175;
wire G398;
wire G172;
wire G51;
wire G421;
wire G490;
wire G510;
wire G341;
wire G373;
wire G213;
wire G465;
wire II493;
wire G444;
wire G354;
wire G344;
wire G300;
wire G47;
wire G320;
wire G57;
wire G488;
wire G239;
wire G419;
wire G414;
wire G312;
wire G227;
wire G392;
wire G162;
wire G197;
wire G164;
wire II624;
wire G66;
wire II692;
wire G359;
wire G364;
wire G404;
wire G499;
wire G141;
wire G123;
wire G56;
wire G343;
wire G268;
wire G97;
wire G271;
wire II386;
wire G435;
wire G150;
wire G379;
wire G474;
wire G225;
wire G135;
wire G60;
wire G82;
wire G290;
wire G188;
wire G84;
wire G303;
wire G397;
wire G240;
wire G470;
wire G247;
wire G89;
wire G257;
wire G442;
wire G212;
wire G98;
wire G55;
wire II316;
wire G443;
wire G372;
wire G183;
wire G511;
wire G500;
wire G48;
wire G336;
wire G173;
wire G452;
wire G108;
wire II502;
wire G449;
wire G479;
wire G180;
wire G323;
wire G543;
wire G100;
wire G521;
wire G52;
wire G124;
wire G120;
wire G299;
wire G368;
wire G207;
wire G273;
wire G515;
wire G487;
wire G524;
wire G258;
wire G129;
wire G492;
wire G193;
wire G160;
wire G184;
wire G256;
wire G132;
wire G380;
wire G424;
wire G158;
wire G436;
wire G113;
wire G272;
wire G403;
wire G319;
wire G222;
wire G486;
wire G189;
wire G219;
wire G441;
wire G338;
wire G115;
wire G480;
wire G417;
wire G374;
wire G243;
wire G544;
wire G157;
wire G512;
wire II276;
wire G67;
wire G107;
wire G437;
wire G496;
wire G402;
wire II295;
wire G90;
wire G501;
wire G279;
wire G262;
wire G277;
wire G215;
wire II287;
wire G223;
wire G362;
wire G75;
wire G396;
wire G292;
wire II330;
wire G235;
wire G142;
wire G352;
wire G346;
wire G461;
wire G288;
wire G206;
wire G304;
wire G101;
wire G121;
wire G469;
wire G523;
wire G261;
wire G159;
wire II573;
wire G255;
wire G321;
wire G259;
wire G531;
wire G68;
wire G311;
wire G185;
wire G337;
wire G192;
wire G195;
wire II371;
wire G330;
wire G204;
wire G168;
wire II327;
wire G318;
wire G422;
wire G328;
wire G59;
wire G274;
wire G357;
wire G477;
wire G394;
wire G226;
wire G224;
wire G99;
wire G460;
wire G116;
wire G112;
wire G411;
wire G448;
wire G287;
wire G459;
wire G306;
wire G534;
wire G182;
wire G170;
wire G214;
wire G76;
wire G133;
wire G242;
wire G440;
wire G345;
wire G513;
wire G401;
wire G194;
wire G232;
wire G497;
wire G514;
wire G278;
wire G491;
wire G143;
wire G305;
wire G355;
wire G429;
wire G472;
wire G106;
wire G178;
wire G333;
wire G50;
wire G381;
wire G167;
wire G430;
wire G291;
wire G361;
wire G462;
wire G234;
wire G138;
wire G438;
wire G541;
wire G217;
wire G200;
wire G456;
wire G254;
wire G353;
wire G77;
wire G93;
wire G191;
wire G105;
wire G144;
wire G329;
wire G147;
wire G493;
wire G297;
wire G117;
wire G506;
wire G447;
wire II631;
wire G485;
wire G176;
wire G210;
wire G457;
wire G284;
wire G325;
wire G526;
wire G221;
wire G400;
wire G307;
wire G386;
wire G554;
wire G187;
wire G118;
wire G130;
wire G54;
wire G478;
wire G348;
wire G87;
wire G69;
wire G426;
wire G533;
wire II536;
wire G314;
wire G126;
wire G517;
wire G366;
wire G377;
wire II156;
wire G169;
wire G111;
wire G171;
wire G263;
wire G385;
wire G233;
wire G450;
wire G324;
wire G507;
wire G166;
wire G525;
wire G446;
wire G216;
wire G282;
wire G471;
wire G439;
wire G286;
wire G369;
wire G145;
wire G253;
wire G136;
wire G494;
wire G464;
wire G332;
wire G391;
wire G190;
wire G245;
wire G155;
wire G128;
wire G409;
wire G308;
wire G285;
wire G420;
wire G431;
wire G94;
wire G91;
wire G423;
wire G316;
wire G104;
wire G458;
wire G360;
wire G484;
wire II576;
wire G384;
wire G205;
wire G536;
wire G92;
wire G375;
wire G376;
wire G201;
wire G264;
wire G416;
wire G294;
wire G276;
wire G63;
wire G527;
wire G339;
wire G509;
wire G78;
wire G553;
wire G127;
wire G156;
wire G252;
wire G110;
wire G88;
wire G425;
wire G475;
wire G119;
wire G131;
wire G516;
wire G331;
wire G347;
wire G418;
wire G70;
wire G363;
wire G495;
wire G413;
wire G95;
wire G315;
wire G463;
wire G79;
wire G244;
wire G445;
wire G351;
wire G427;
wire G236;
wire G393;
wire G248;
wire G137;
wire G165;
wire G538;
wire G529;
wire G383;
wire G483;
wire G432;
wire G504;
wire G174;
wire G342;
wire G146;
wire G309;
wire G378;
wire G198;
wire G289;
wire G408;
wire G387;
wire G73;
wire G163;
wire G251;
wire G148;
wire G153;
wire G85;
wire G519;
wire G74;
wire G230;
wire G283;
wire G103;
wire G326;
wire G49;
wire G177;
wire II529;
wire G208;
wire G211;
wire G293;
wire G265;
wire G71;
wire G410;
wire G267;
wire G275;
wire G406;
wire G520;
wire G335;
wire G281;
wire G322;
wire G202;
wire G358;
wire II374;
wire G508;
wire G370;
wire G149;
wire G468;
wire G139;
wire G109;
wire G237;
wire G528;
wire G428;
wire II249;
wire G473;
wire G125;
wire G181;
wire G298;
wire G454;
wire G476;
wire G350;
wire G229;
wire G296;
wire G199;
wire G399;
wire G482;
wire II272;
wire G179;
wire G62;
wire G102;
wire G502;
wire G317;
wire G152;
wire II352;
wire G382;
wire G388;
wire G64;
wire G250;
wire G86;
wire G241;
wire G334;
wire G505;
wire G407;
wire G231;
wire G280;
wire G415;
wire G327;
wire G72;
wire G266;
wire G203;
wire G455;
wire G186;
wire G96;
wire G53;
wire G451;
wire G249;
wire II280;
wire II662;
wire G220;
wire G540;
wire G390;
wire G367;
wire G349;
wire G433;
wire G545;
wire G518;
wire G340;
wire G154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G29 <= 0;
  else
    G29 <= G502;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G30 <= 0;
  else
    G30 <= G503;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G31 <= 0;
  else
    G31 <= G504;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G32 <= 0;
  else
    G32 <= G505;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G33 <= 0;
  else
    G33 <= G506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G34 <= 0;
  else
    G34 <= G507;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G35 <= 0;
  else
    G35 <= G508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G36 <= 0;
  else
    G36 <= G509;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G37 <= 0;
  else
    G37 <= G510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G38 <= 0;
  else
    G38 <= G511;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G39 <= 0;
  else
    G39 <= G512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G40 <= 0;
  else
    G40 <= G513;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G41 <= 0;
  else
    G41 <= G514;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G42 <= 0;
  else
    G42 <= G515;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G43 <= 0;
  else
    G43 <= G516;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G44 <= 0;
  else
    G44 <= G517;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G45 <= 0;
  else
    G45 <= G518;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    G46 <= 0;
  else
    G46 <= G519;
assign G260 = ((~G528))|((~G529))|((~G191));
assign G228 = ((~G524));
assign G196 = ((~G5)&(~G540)&(~G86));
assign G61 = (G405)|(G406);
assign G546 = ((~G41));
assign G140 = ((~G33));
assign G371 = (G161&G168&G267);
assign G489 = ((~G273));
assign G498 = ((~G195));
assign G161 = ((~G316))|((~G72));
assign G301 = (G122)|(G486);
assign G395 = (G4)|(G134);
assign G453 = (G545&G186);
assign G209 = ((~G1)&(~G524));
assign G365 = (G282&G137&G156);
assign G356 = (G6)|(G476);
assign G295 = (G122)|(G491);
assign G313 = (G521)|(G475);
assign G270 = ((~G345))|((~G204));
assign G522 = ((~G2));
assign G218 = ((~G528)&(~G217));
assign G134 = ((~G3))|((~G5));
assign G269 = (G362)|(G529);
assign G83 = ((~G355))|((~G356));
assign G80 = ((~G421))|((~G226))|((~G256));
assign G122 = ((~G522))|((~G3));
assign G503 = ((~G286))|((~G538));
assign G389 = (G9)|(G274);
assign G151 = ((~G305))|((~G200));
assign G412 = (G3&G207);
assign G405 = ((~II662));
assign G81 = (G288&G240);
assign G58 = ((~G1))|((~G3));
assign G434 = (G165&G231);
assign G310 = (G522)|(G135);
assign G238 = ((~G2))|((~G524));
assign G114 = (G385)|(G386);
assign II218 = ((~G528));
assign G302 = (G4)|(G529);
assign G246 = ((~G544))|((~G186));
assign G175 = ((~G86)&(~G500));
assign G398 = (G94&G156&G158);
assign G172 = ((~G171));
assign G51 = ((~G260))|((~G237));
assign G421 = (G521)|(G2)|(G228);
assign G490 = ((~G190));
assign G510 = ((~G350))|((~G235));
assign G341 = (G531&G118);
assign G373 = (G34&G160);
assign G213 = ((~G64))|((~G275));
assign G465 = (G524)|(G210);
assign II493 = ((~G218));
assign G444 = (G64&G78&G211);
assign G354 = (G0&G214);
assign G344 = (G111&G189&G195);
assign G300 = (G87)|(G97);
assign G47 = (G440)|(G441);
assign G320 = (G76)|(G272);
assign G57 = ((~G0))|((~G2));
assign G488 = ((~G172));
assign G239 = ((~G7))|((~G533));
assign G419 = (G3)|(G5);
assign G312 = (G180&G182);
assign G414 = ((~II386));
assign G227 = ((~G5)&(~G200));
assign G551 = (G327)|(G328)|(G329);
assign G392 = (G132&G155);
assign G539 = (G451)|(G452)|(G453);
assign G162 = ((~G185)&(~G498));
assign G197 = ((~G540)&(~G232));
assign G164 = ((~G531)&(~G10));
assign II624 = ((~G120));
assign G66 = ((~G129))|((~G101));
assign II692 = ((~G145));
assign G359 = (G6&G31);
assign G364 = (G2&G109);
assign G404 = ((~II493));
assign G141 = (G353)|(G354);
assign G499 = ((~G280));
assign G123 = ((~G122));
assign G56 = ((~G374))|((~G375));
assign G343 = (G2&G528&G147);
assign G268 = ((~G11))|((~G113));
assign G97 = ((~G2))|((~G5));
assign G271 = ((~G1))|((~G4));
assign II386 = ((~G199));
assign G435 = ((~II327));
assign G150 = (G303)|(G304);
assign G379 = (G9&G211);
assign G474 = (G242&G77);
assign G225 = ((~G7)&(~G8));
assign G135 = ((~G134));
assign G60 = (G413)|(G414);
assign G82 = ((~G334))|((~G335));
assign G290 = (G117&G135&G157);
assign G188 = ((~G543)&(~G493));
assign G84 = ((~G369))|((~G370));
assign G303 = ((~II624));
assign G397 = (G101&G98&G157);
assign G240 = ((~G4))|((~G134));
assign G470 = (G528&G149);
assign G247 = ((~G471)&(~G472)&(~G473)&(~G474));
assign G89 = ((~G531))|((~G8));
assign G257 = ((~G538))|((~G230));
assign G442 = (G541&G121);
assign G212 = ((~G213));
assign G98 = ((~G97));
assign G55 = ((~G54));
assign II316 = ((~G239));
assign G443 = (G47&G162);
assign G372 = (G116&G275&G155);
assign G183 = ((~G330)&(~G3));
assign G511 = (G163&G164);
assign G500 = ((~G173));
assign G532 = (G422)|(G423);
assign G48 = ((~G407))|((~G408))|((~G409));
assign G452 = (G526&G184);
assign G336 = ((~II631));
assign G173 = ((~G495));
assign G108 = (G346)|(G347);
assign II502 = ((~G124));
assign G449 = (G88&G154);
assign G479 = ((~G194));
assign G180 = ((~G181));
assign G323 = (G2&G144);
assign G543 = ((~G13));
assign G100 = ((~G381))|((~G220));
assign G521 = ((~G1));
assign G52 = ((~G298))|((~G299))|((~G219));
assign G124 = ((~G206));
assign G120 = ((~G294))|((~G295));
assign G299 = ((~II352));
assign G368 = (G533)|(G536);
assign G207 = ((~G208));
assign G273 = ((~G325))|((~G326));
assign G515 = ((~G387)&(~G388));
assign G487 = ((~G534));
assign G524 = ((~G3));
assign G258 = ((~G464))|((~G103))|((~G223));
assign G129 = ((~G527))|((~G5));
assign G492 = ((~G62));
assign G193 = (G6)|(G30);
assign G160 = ((~G161));
assign G184 = ((~G541)&(~G13)&(~G499));
assign G256 = ((~G4))|((~G69));
assign G132 = ((~G42));
assign G380 = (G6&G93);
assign G424 = (G78&G174&G177);
assign G158 = ((~G521)&(~G281));
assign G436 = (G123&G77);
assign G113 = ((~G389))|((~G390));
assign G272 = ((~G271));
assign G403 = ((~II573));
assign G319 = (G529)|(G489);
assign G222 = ((~G533))|((~G10));
assign G486 = ((~G68));
assign G189 = ((~G522)&(~G54));
assign G219 = ((~G524))|((~G55));
assign G441 = ((~II330));
assign G338 = (G202&G203);
assign G115 = (G457)|(G458)|(G459);
assign G480 = ((~G179));
assign G417 = (G13&G282&G70);
assign G243 = ((~G368))|((~G275))|((~G34));
assign G374 = (G536)|(G538);
assign G544 = (G343)|(G344);
assign G157 = ((~G13)&(~G483));
assign G512 = ((~G310))|((~G233));
assign II276 = ((~G238));
assign G67 = ((~G44));
assign G107 = ((~G456));
assign G437 = (G66&G229);
assign G549 = (G396)|(G397)|(G398)|(G477);
assign G402 = (G154&G183);
assign G496 = ((~G188));
assign II295 = ((~G198));
assign G90 = ((~G89));
assign G501 = ((~G156));
assign G279 = (G317)|(G166);
assign G262 = ((~G527))|((~G278));
assign G277 = ((~G394))|((~G395))|((~G81));
assign G215 = ((~G135))|((~G55))|((~G212));
assign II287 = ((~G135));
assign G223 = ((~G224));
assign G362 = (G129&G77);
assign G75 = ((~G74));
assign G396 = (G76&G272&G155);
assign G292 = (G538)|(G75);
assign II330 = ((~G236));
assign G235 = ((~G6))|((~G536));
assign G142 = (G403)|(G404);
assign G352 = (G8&G135&G37&G164);
assign G346 = (G2&G82);
assign G461 = (G529&G531);
assign G206 = ((~G287))|((~G524));
assign G288 = (G1)|(G528);
assign G304 = (G52&G158);
assign G101 = ((~G3))|((~G4));
assign G121 = (G438)|(G439);
assign G523 = ((~G254))|((~G255))|((~G208));
assign G469 = (G163&G3);
assign G261 = (G283)|(G528);
assign G159 = ((~G6))|((~G155));
assign II573 = ((~G176));
assign G255 = ((~G309))|((~G2))|((~G529));
assign G321 = (G90&G50);
assign G259 = ((~G130))|((~G225));
assign G531 = ((~G7));
assign G68 = ((~G302))|((~G528));
assign G185 = ((~G525))|((~G184));
assign G311 = (G0&G178&G179);
assign G337 = (G270&G167);
assign G192 = ((~G193));
assign G195 = ((~G521)&(~G134));
assign II371 = ((~G1));
assign G330 = (G248&G249);
assign G204 = ((~G521))|((~G87));
assign II327 = ((~G135));
assign G168 = ((~G75))|((~G221));
assign G318 = (G6)|(G8)|(G232);
assign G422 = (G0&G80&G155);
assign G328 = (G5&G102&G155);
assign G59 = ((~G58));
assign G274 = ((~G7))|((~G10));
assign G477 = ((~G276));
assign G357 = (G265&G232);
assign G394 = (G5)|(G58);
assign G226 = ((~G527))|((~G59));
assign G224 = (G533)|(G31);
assign G99 = ((~G29));
assign G460 = (G2&G81&G115);
assign G116 = ((~G6))|((~G9));
assign G112 = ((~G8))|((~G31));
assign G411 = (G48&G59);
assign G448 = (G139&G153);
assign G287 = (G522)|(G81);
assign G459 = ((~II295));
assign G306 = (G524&G78);
assign G534 = ((~G296))|((~G297))|((~G166));
assign G182 = ((~G12)&(~G62));
assign G170 = ((~G171));
assign G214 = ((~G215));
assign G76 = ((~G0))|((~G3));
assign G133 = (G434)|(G435);
assign G242 = (G469)|(G470);
assign G440 = (G38&G234);
assign G345 = (G529)|(G226);
assign G550 = (G289)|(G290)|(G291)|(G485);
assign G513 = ((~G360)&(~G361));
assign G401 = (G2&G110&G155);
assign G232 = ((~G536))|((~G164));
assign G194 = ((~G281)&(~G271));
assign G497 = ((~G205));
assign G514 = ((~G372)&(~G373)&(~G478));
assign G278 = ((~G332))|((~G333));
assign G491 = ((~G194));
assign G305 = (G524)|(G55);
assign G143 = ((~G258))|((~G193))|((~G259));
assign G355 = (G11)|(G116);
assign G429 = (G51&G225);
assign G472 = (G136&G9&G190);
assign G106 = (G358)|(G359);
assign G178 = ((~G521)&(~G4));
assign G333 = ((~II218));
assign G50 = ((~G49));
assign G381 = (G7)|(G71);
assign G167 = ((~G168));
assign G430 = (G177&G196);
assign G234 = ((~G235));
assign G462 = (G192&G538);
assign G361 = (G6&G202);
assign G291 = (G138&G155);
assign G138 = ((~G465))|((~G263));
assign G438 = (G8&G146&G133);
assign G541 = ((~G12));
assign G217 = ((~G50))|((~G230));
assign G200 = ((~G527))|((~G529));
assign G456 = ((~II374));
assign G254 = ((~G1))|((~G152));
assign G353 = (G11&G92&G163);
assign G77 = ((~G4))|((~G528));
assign G93 = (G376)|(G377)|(G378);
assign G191 = ((~G9)&(~G482));
assign G105 = (G321)|(G273);
assign G144 = ((~G215))|((~G252))|((~G253));
assign G329 = (G150&G156);
assign G147 = (G341)|(G342);
assign G493 = ((~G544));
assign G297 = (G64)|(G274);
assign G117 = ((~G2))|((~G4));
assign G506 = ((~G311)&(~G312));
assign G447 = ((~II576));
assign II631 = ((~G188));
assign G485 = ((~G276));
assign G176 = ((~G4)&(~G494));
assign G210 = ((~G520))|((~G272));
assign G457 = (G4&G107);
assign G284 = (G528)|(G272)|(G281);
assign G526 = ((~G1))|((~G2))|((~G141));
assign G325 = (G7)|(G536)|(G222);
assign G221 = ((~G222));
assign G400 = (G0&G277);
assign G307 = (G6&G104);
assign G386 = (G536&G85);
assign G554 = ((~G553));
assign G187 = ((~G13)&(~G492));
assign G118 = (G337)|(G338);
assign G130 = ((~G9));
assign G54 = ((~G4))|((~G6));
assign G478 = ((~G279));
assign G348 = (G97&G55);
assign G87 = ((~G86));
assign G69 = ((~G419))|((~G420))|((~G233));
assign G426 = (G37&G162&G38);
assign G533 = ((~G8));
assign II536 = ((~G79));
assign G126 = (G363)|(G364);
assign G314 = (G527)|(G57);
assign G517 = ((~G428)&(~G429));
assign G366 = (G125&G155);
assign G377 = (G90&G56);
assign II156 = ((~G4));
assign G169 = ((~G5)&(~G7));
assign G111 = ((~G213))|((~G217));
assign G171 = ((~G553))|((~G187));
assign G263 = ((~G0))|((~G99));
assign G385 = (G529&G7&G49);
assign G233 = ((~G522))|((~G135));
assign G450 = (G12)|(G171);
assign G324 = (G522&G183);
assign G507 = ((~G315)&(~G12)&(~G487));
assign G166 = ((~G7))|((~G50));
assign G525 = ((~G526));
assign G446 = ((~II536));
assign G216 = ((~G4)&(~G5));
assign G282 = ((~G281));
assign G471 = (G191&G103&G112);
assign G439 = (G174&G175);
assign G286 = (G9)|(G540);
assign G369 = ((~II316));
assign G253 = ((~G87))|((~G218));
assign G145 = (G426)|(G427);
assign G136 = ((~G222))|((~G224));
assign G494 = ((~G173));
assign G464 = (G72)|(G536);
assign G332 = ((~II276));
assign G391 = (G74)|(G220);
assign G190 = ((~G7)&(~G11));
assign G155 = ((~G13)&(~G480));
assign G245 = ((~G8))|((~G34));
assign G128 = (G415)|(G416)|(G417)|(G418);
assign G409 = (G528)|(G55);
assign G308 = (G5&G151);
assign G285 = (G5)|(G479);
assign G431 = (G524&G67);
assign G420 = (G522)|(G59);
assign G94 = ((~G261))|((~G181))|((~G262));
assign G91 = (G430)|(G431);
assign G423 = (G541&G128);
assign G542 = ((~G243))|((~G244))|((~G279));
assign G104 = ((~G122))|((~G238))|((~G240));
assign G316 = (G531)|(G536);
assign G458 = ((~II272));
assign G360 = (G8&G106);
assign G484 = ((~G30));
assign II576 = ((~G175));
assign G384 = (G529)|(G71);
assign G205 = ((~G529)&(~G122));
assign G536 = ((~G9));
assign G92 = (G351)|(G352);
assign G375 = (G10)|(G540);
assign G376 = (G533&G75);
assign G201 = ((~G528)&(~G54));
assign G264 = ((~G227))|((~G241));
assign G416 = (G61&G167);
assign G294 = (G1)|(G117)|(G281);
assign G276 = ((~G3))|((~G543))|((~G140));
assign G63 = ((~G75))|((~G8));
assign G527 = ((~G4));
assign G339 = (G533&G199&G209);
assign G509 = ((~G331)&(~G5));
assign G78 = ((~G77));
assign G547 = (G382)|(G383);
assign G553 = (G322)|(G323)|(G324);
assign G127 = ((~G391))|((~G268));
assign G156 = ((~G12)&(~G543));
assign G252 = ((~G3))|((~G11))|((~G35))|((~G216));
assign G110 = (G399)|(G400);
assign G88 = (G446)|(G447);
assign G425 = (G146&G176);
assign G475 = ((~G57));
assign G119 = ((~G284))|((~G285));
assign G131 = (G379)|(G380);
assign G516 = ((~G410)&(~G411)&(~G412));
assign G331 = (G213&G257);
assign G347 = ((~II287));
assign G418 = (G524&G60&G172);
assign G70 = ((~G43));
assign G363 = (G77&G205);
assign G495 = ((~G273));
assign G413 = (G197&G201);
assign G95 = (G424)|(G425);
assign G552 = (G365)|(G366)|(G367);
assign G315 = (G250&G251);
assign G463 = (G521&G148);
assign G79 = (G444)|(G445);
assign G244 = (G371)|(G159);
assign G445 = (G53&G225);
assign G351 = (G524&G169&G221&G234);
assign G427 = (G541&G95&G165);
assign G236 = ((~G274));
assign G393 = (G127&G34);
assign G248 = ((~G529))|((~G36));
assign G137 = (G348)|(G349);
assign G165 = ((~G529));
assign G538 = ((~G10));
assign G529 = ((~G6));
assign G383 = (G131&G155);
assign G483 = ((~G182));
assign G432 = ((~II692));
assign G504 = ((~G292))|((~G293));
assign G174 = ((~G496));
assign G342 = (G73&G197);
assign G309 = ((~II280));
assign G378 = (G89&G50);
assign G146 = (G336)|(G170);
assign G198 = ((~G520)&(~G3));
assign G289 = (G2&G119&G156);
assign G408 = (G529)|(G77);
assign G387 = (G6&G274&G75);
assign G73 = (G339)|(G340);
assign G163 = ((~G0)&(~G4));
assign G251 = ((~G543))|((~G32));
assign G148 = ((~G454))|((~G455))|((~G0));
assign G153 = ((~G522));
assign G85 = ((~G384))|((~G239));
assign G519 = ((~G460)&(~G461)&(~G462)&(~G463));
assign G230 = ((~G8)&(~G490));
assign G74 = ((~G9))|((~G11));
assign G283 = (G122&G219);
assign G103 = ((~G529))|((~G7))|((~G30));
assign G326 = (G533)|(G232);
assign G49 = ((~G9))|((~G538));
assign II529 = ((~G468));
assign G177 = ((~G357));
assign G208 = ((~G68))|((~G229));
assign G211 = ((~G6)&(~G274));
assign G548 = (G392)|(G393);
assign G293 = (G7)|(G540);
assign G265 = ((~G50));
assign G410 = (G1&G205);
assign G71 = ((~G8))|((~G10));
assign G267 = ((~G536))|((~G84));
assign G275 = ((~G274));
assign G406 = (G87&G172);
assign G520 = ((~G0));
assign G335 = ((~II371));
assign G281 = ((~G523))|((~G534));
assign G322 = (G522&G105&G196);
assign G202 = ((~G10)&(~G63));
assign G358 = (G7&G83);
assign II374 = ((~G520));
assign G508 = ((~G318))|((~G319));
assign G535 = (G432)|(G433);
assign G370 = ((~II249));
assign G149 = ((~II529));
assign G468 = ((~II502));
assign G139 = (G442)|(G443);
assign G109 = ((~G269))|((~G219));
assign G537 = (G448)|(G449);
assign G237 = ((~G10))|((~G75))|((~G201));
assign G528 = ((~G5));
assign G428 = (G212&G227);
assign II249 = ((~G538));
assign G473 = (G11&G143);
assign G125 = ((~G40));
assign G181 = ((~G2))|((~G78));
assign G298 = (G5)|(G497);
assign G454 = (G122)|(G77);
assign G476 = ((~G30));
assign G350 = (G6)|(G536);
assign G229 = ((~G1)&(~G522));
assign G296 = (G89)|(G484);
assign G199 = ((~G200));
assign G399 = (G520&G1);
assign G482 = ((~G241));
assign G179 = ((~G541)&(~G280));
assign II272 = ((~G209));
assign G62 = ((~G534))|((~G32));
assign G502 = ((~G436)&(~G437));
assign G102 = ((~G320))|((~G266))|((~G210));
assign G317 = (G159&G245);
assign II352 = ((~G77));
assign G382 = (G9&G100&G34);
assign G388 = (G11&G114);
assign G152 = (G306)|(G307)|(G308);
assign G64 = ((~G63));
assign G250 = ((~G13))|((~G523));
assign G86 = ((~G55))|((~G3));
assign G241 = ((~G10)&(~G11));
assign G334 = ((~II156));
assign G505 = ((~G300))|((~G301))|((~G181));
assign G407 = (G6)|(G117);
assign G231 = ((~G232));
assign G280 = ((~G46))|((~G247));
assign G415 = (G146&G142&G165);
assign G327 = (G4&G39&G157);
assign G72 = ((~G71));
assign G266 = ((~G524))|((~G96));
assign G203 = ((~G204));
assign G186 = ((~G282)&(~G501));
assign G455 = (G78)|(G206);
assign G96 = ((~G313))|((~G314));
assign G53 = ((~G264))|((~G237));
assign G451 = (G541&G554&G187);
assign G249 = ((~G11))|((~G273))|((~G201));
assign II280 = ((~G272));
assign II662 = ((~G174));
assign G220 = ((~G7))|((~G71));
assign G540 = ((~G11));
assign G390 = (G89)|(G50);
assign G367 = (G126&G157);
assign G349 = (G6&G108);
assign G433 = (G91&G154);
assign G545 = ((~G544));
assign G530 = (G401)|(G402);
assign G518 = ((~G450))|((~G185))|((~G246));
assign G340 = (G8&G270);
assign G154 = ((~G12)&(~G488));
endmodule
