module s38417(
  blif_clk_net,
  blif_reset_net,
  g51,
  g563,
  g1249,
  g1943,
  g2637,
  g3212,
  g3213,
  g3214,
  g3215,
  g3216,
  g3217,
  g3218,
  g3219,
  g3220,
  g3221,
  g3222,
  g3223,
  g3224,
  g3225,
  g3226,
  g3227,
  g3228,
  g3229,
  g3230,
  g3231,
  g3232,
  g3233,
  g3234,
  g3993,
  g4088,
  g4090,
  g4200,
  g4321,
  g4323,
  g4450,
  g4590,
  g5388,
  g5437,
  g5472,
  g5511,
  g5549,
  g5555,
  g5595,
  g5612,
  g5629,
  g5637,
  g5648,
  g5657,
  g5686,
  g5695,
  g5738,
  g5747,
  g5796,
  g6225,
  g6231,
  g6313,
  g6368,
  g6442,
  g6447,
  g6485,
  g6518,
  g6573,
  g6642,
  g6677,
  g6712,
  g6750,
  g6782,
  g6837,
  g6895,
  g6911,
  g6944,
  g6979,
  g7014,
  g7052,
  g7084,
  g7161,
  g7194,
  g7229,
  g7264,
  g7302,
  g7334,
  g7357,
  g7390,
  g7425,
  g7487,
  g7519,
  g7909,
  g7956,
  g7961,
  g8007,
  g8012,
  g8021,
  g8023,
  g8030,
  g8082,
  g8087,
  g8096,
  g8106,
  g8167,
  g8175,
  g8249,
  g8251,
  g8258,
  g8259,
  g8260,
  g8261,
  g8262,
  g8263,
  g8264,
  g8265,
  g8266,
  g8267,
  g8268,
  g8269,
  g8270,
  g8271,
  g8272,
  g8273,
  g8274,
  g8275,
  g16297,
  g16355,
  g16399,
  g16437,
  g16496,
  g24734,
  g25420,
  g25435,
  g25442,
  g25489,
  g26104,
  g26135,
  g26149,
  g27380);
input blif_clk_net;
input blif_reset_net;
input g51;
input g563;
input g1249;
input g1943;
input g2637;
input g3212;
input g3213;
input g3214;
input g3215;
input g3216;
input g3217;
input g3218;
input g3219;
input g3220;
input g3221;
input g3222;
input g3223;
input g3224;
input g3225;
input g3226;
input g3227;
input g3228;
input g3229;
input g3230;
input g3231;
input g3232;
input g3233;
input g3234;
output g3993;
output g4088;
output g4090;
output g4200;
output g4321;
output g4323;
output g4450;
output g4590;
output g5388;
output g5437;
output g5472;
output g5511;
output g5549;
output g5555;
output g5595;
output g5612;
output g5629;
output g5637;
output g5648;
output g5657;
output g5686;
output g5695;
output g5738;
output g5747;
output g5796;
output g6225;
output g6231;
output g6313;
output g6368;
output g6442;
output g6447;
output g6485;
output g6518;
output g6573;
output g6642;
output g6677;
output g6712;
output g6750;
output g6782;
output g6837;
output g6895;
output g6911;
output g6944;
output g6979;
output g7014;
output g7052;
output g7084;
output g7161;
output g7194;
output g7229;
output g7264;
output g7302;
output g7334;
output g7357;
output g7390;
output g7425;
output g7487;
output g7519;
output g7909;
output g7956;
output g7961;
output g8007;
output g8012;
output g8021;
output g8023;
output g8030;
output g8082;
output g8087;
output g8096;
output g8106;
output g8167;
output g8175;
output g8249;
output g8251;
output g8258;
output g8259;
output g8260;
output g8261;
output g8262;
output g8263;
output g8264;
output g8265;
output g8266;
output g8267;
output g8268;
output g8269;
output g8270;
output g8271;
output g8272;
output g8273;
output g8274;
output g8275;
output g16297;
output g16355;
output g16399;
output g16437;
output g16496;
output g24734;
output g25420;
output g25435;
output g25442;
output g25489;
output g26104;
output g26135;
output g26149;
output g27380;
reg g2814;
reg g2817;
reg g2933;
reg g2950;
reg g2883;
reg g2888;
reg g2896;
reg g2892;
reg g2903;
reg g2900;
reg g2908;
reg g2912;
reg g2917;
reg g2924;
reg g2920;
reg g2984;
reg g2985;
reg g2930;
reg g2929;
reg g2879;
reg g2934;
reg g2935;
reg g2938;
reg g2941;
reg g2944;
reg g2947;
reg g2953;
reg g2956;
reg g2959;
reg g2962;
reg g2963;
reg g2966;
reg g2969;
reg g2972;
reg g2975;
reg g2978;
reg g2981;
reg g2874;
reg g1506;
reg g1501;
reg g1496;
reg g1491;
reg g1486;
reg g1481;
reg g1476;
reg g1471;
reg g2877;
reg g2861;
reg g813;
reg g2864;
reg g809;
reg g2867;
reg g805;
reg g2870;
reg g801;
reg g2818;
reg g797;
reg g2821;
reg g793;
reg g2824;
reg g789;
reg g2827;
reg g785;
reg g2830;
reg g2873;
reg g2833;
reg g125;
reg g2836;
reg g121;
reg g2839;
reg g117;
reg g2842;
reg g113;
reg g2845;
reg g109;
reg g2848;
reg g105;
reg g2851;
reg g101;
reg g2854;
reg g97;
reg g2858;
reg g2857;
reg g2200;
reg g2195;
reg g2190;
reg g2185;
reg g2180;
reg g2175;
reg g2170;
reg g2165;
reg g2878;
reg g3129;
reg g3117;
reg g3109;
reg g3210;
reg g3211;
reg g3084;
reg g3085;
reg g3086;
reg g3087;
reg g3091;
reg g3092;
reg g3093;
reg g3094;
reg g3095;
reg g3096;
reg g3097;
reg g3098;
reg g3099;
reg g3100;
reg g3101;
reg g3102;
reg g3103;
reg g3104;
reg g3105;
reg g3106;
reg g3107;
reg g3108;
reg g3155;
reg g3158;
reg g3161;
reg g3164;
reg g3167;
reg g3170;
reg g3173;
reg g3176;
reg g3179;
reg g3182;
reg g3185;
reg g3088;
reg g3191;
reg g3194;
reg g3197;
reg g3198;
reg g3201;
reg g3204;
reg g3207;
reg g3188;
reg g3133;
reg g3132;
reg g3128;
reg g3127;
reg g3126;
reg g3125;
reg g3124;
reg g3123;
reg g3120;
reg g3114;
reg g3113;
reg g3112;
reg g3110;
reg g3111;
reg g3139;
reg g3136;
reg g3134;
reg g3135;
reg g3151;
reg g3142;
reg g3147;
reg g185;
reg g138;
reg g135;
reg g165;
reg g130;
reg g131;
reg g129;
reg g133;
reg g134;
reg g132;
reg g142;
reg g143;
reg g141;
reg g145;
reg g146;
reg g144;
reg g148;
reg g149;
reg g147;
reg g151;
reg g152;
reg g150;
reg g154;
reg g155;
reg g153;
reg g157;
reg g158;
reg g156;
reg g160;
reg g161;
reg g159;
reg g163;
reg g164;
reg g162;
reg g169;
reg g170;
reg g168;
reg g172;
reg g173;
reg g171;
reg g175;
reg g176;
reg g174;
reg g178;
reg g179;
reg g177;
reg g186;
reg g189;
reg g192;
reg g231;
reg g234;
reg g237;
reg g195;
reg g198;
reg g201;
reg g240;
reg g243;
reg g246;
reg g204;
reg g207;
reg g210;
reg g249;
reg g252;
reg g255;
reg g213;
reg g216;
reg g219;
reg g258;
reg g261;
reg g264;
reg g222;
reg g225;
reg g228;
reg g267;
reg g270;
reg g273;
reg g92;
reg g88;
reg g83;
reg g79;
reg g74;
reg g70;
reg g65;
reg g61;
reg g56;
reg g52;
reg g180;
reg g182;
reg g181;
reg g276;
reg g405;
reg g401;
reg g309;
reg g354;
reg g343;
reg g346;
reg g369;
reg g358;
reg g361;
reg g384;
reg g373;
reg g376;
reg g398;
reg g388;
reg g391;
reg g408;
reg g411;
reg g414;
reg g417;
reg g420;
reg g423;
reg g427;
reg g428;
reg g426;
reg g429;
reg g432;
reg g435;
reg g438;
reg g441;
reg g444;
reg g448;
reg g449;
reg g447;
reg g312;
reg g313;
reg g314;
reg g315;
reg g316;
reg g317;
reg g318;
reg g319;
reg g320;
reg g322;
reg g323;
reg g321;
reg g403;
reg g404;
reg g402;
reg g450;
reg g451;
reg g452;
reg g453;
reg g454;
reg g279;
reg g280;
reg g281;
reg g282;
reg g283;
reg g284;
reg g285;
reg g286;
reg g287;
reg g288;
reg g289;
reg g290;
reg g291;
reg g299;
reg g305;
reg g308;
reg g297;
reg g296;
reg g295;
reg g294;
reg g304;
reg g303;
reg g302;
reg g301;
reg g300;
reg g298;
reg g342;
reg g349;
reg g350;
reg g351;
reg g352;
reg g353;
reg g357;
reg g364;
reg g365;
reg g366;
reg g367;
reg g368;
reg g372;
reg g379;
reg g380;
reg g381;
reg g382;
reg g383;
reg g387;
reg g394;
reg g395;
reg g396;
reg g397;
reg g324;
reg g325;
reg g331;
reg g337;
reg g545;
reg g551;
reg g550;
reg g554;
reg g557;
reg g510;
reg g513;
reg g523;
reg g524;
reg g564;
reg g569;
reg g570;
reg g571;
reg g572;
reg g573;
reg g574;
reg g565;
reg g566;
reg g567;
reg g568;
reg g489;
reg g474;
reg g481;
reg g485;
reg g486;
reg g487;
reg g488;
reg g455;
reg g458;
reg g461;
reg g477;
reg g478;
reg g479;
reg g480;
reg g484;
reg g464;
reg g465;
reg g468;
reg g471;
reg g528;
reg g535;
reg g542;
reg g543;
reg g544;
reg g548;
reg g549;
reg g499;
reg g558;
reg g559;
reg g576;
reg g577;
reg g575;
reg g579;
reg g580;
reg g578;
reg g582;
reg g583;
reg g581;
reg g585;
reg g586;
reg g584;
reg g587;
reg g590;
reg g593;
reg g596;
reg g599;
reg g602;
reg g614;
reg g617;
reg g620;
reg g605;
reg g608;
reg g611;
reg g490;
reg g493;
reg g496;
reg g506;
reg g507;
reg g508;
reg g509;
reg g514;
reg g515;
reg g516;
reg g517;
reg g518;
reg g519;
reg g520;
reg g525;
reg g529;
reg g530;
reg g531;
reg g532;
reg g533;
reg g534;
reg g536;
reg g537;
reg g538;
reg g541;
reg g623;
reg g626;
reg g629;
reg g630;
reg g659;
reg g640;
reg g633;
reg g653;
reg g646;
reg g660;
reg g672;
reg g666;
reg g679;
reg g686;
reg g692;
reg g699;
reg g700;
reg g698;
reg g702;
reg g703;
reg g701;
reg g705;
reg g706;
reg g704;
reg g708;
reg g709;
reg g707;
reg g711;
reg g712;
reg g710;
reg g714;
reg g715;
reg g713;
reg g717;
reg g718;
reg g716;
reg g720;
reg g721;
reg g719;
reg g723;
reg g724;
reg g722;
reg g726;
reg g727;
reg g725;
reg g729;
reg g730;
reg g728;
reg g732;
reg g733;
reg g731;
reg g735;
reg g736;
reg g734;
reg g738;
reg g739;
reg g737;
reg g826;
reg g823;
reg g853;
reg g818;
reg g819;
reg g817;
reg g821;
reg g822;
reg g820;
reg g830;
reg g831;
reg g829;
reg g833;
reg g834;
reg g832;
reg g836;
reg g837;
reg g835;
reg g839;
reg g840;
reg g838;
reg g842;
reg g843;
reg g841;
reg g845;
reg g846;
reg g844;
reg g848;
reg g849;
reg g847;
reg g851;
reg g852;
reg g850;
reg g857;
reg g858;
reg g856;
reg g860;
reg g861;
reg g859;
reg g863;
reg g864;
reg g862;
reg g866;
reg g867;
reg g865;
reg g873;
reg g876;
reg g879;
reg g918;
reg g921;
reg g924;
reg g882;
reg g885;
reg g888;
reg g927;
reg g930;
reg g933;
reg g891;
reg g894;
reg g897;
reg g936;
reg g939;
reg g942;
reg g900;
reg g903;
reg g906;
reg g945;
reg g948;
reg g951;
reg g909;
reg g912;
reg g915;
reg g954;
reg g957;
reg g960;
reg g780;
reg g776;
reg g771;
reg g767;
reg g762;
reg g758;
reg g753;
reg g749;
reg g744;
reg g740;
reg g868;
reg g870;
reg g869;
reg g963;
reg g1092;
reg g1088;
reg g996;
reg g1041;
reg g1030;
reg g1033;
reg g1056;
reg g1045;
reg g1048;
reg g1071;
reg g1060;
reg g1063;
reg g1085;
reg g1075;
reg g1078;
reg g1095;
reg g1098;
reg g1101;
reg g1104;
reg g1107;
reg g1110;
reg g1114;
reg g1115;
reg g1113;
reg g1116;
reg g1119;
reg g1122;
reg g1125;
reg g1128;
reg g1131;
reg g1135;
reg g1136;
reg g1134;
reg g999;
reg g1000;
reg g1001;
reg g1002;
reg g1003;
reg g1004;
reg g1005;
reg g1006;
reg g1007;
reg g1009;
reg g1010;
reg g1008;
reg g1090;
reg g1091;
reg g1089;
reg g1137;
reg g1138;
reg g1139;
reg g1140;
reg g1141;
reg g966;
reg g967;
reg g968;
reg g969;
reg g970;
reg g971;
reg g972;
reg g973;
reg g974;
reg g975;
reg g976;
reg g977;
reg g978;
reg g986;
reg g992;
reg g995;
reg g984;
reg g983;
reg g982;
reg g981;
reg g991;
reg g990;
reg g989;
reg g988;
reg g987;
reg g985;
reg g1029;
reg g1036;
reg g1037;
reg g1038;
reg g1039;
reg g1040;
reg g1044;
reg g1051;
reg g1052;
reg g1053;
reg g1054;
reg g1055;
reg g1059;
reg g1066;
reg g1067;
reg g1068;
reg g1069;
reg g1070;
reg g1074;
reg g1081;
reg g1082;
reg g1083;
reg g1084;
reg g1011;
reg g1012;
reg g1018;
reg g1024;
reg g1231;
reg g1237;
reg g1236;
reg g1240;
reg g1243;
reg g1196;
reg g1199;
reg g1209;
reg g1210;
reg g1250;
reg g1255;
reg g1256;
reg g1257;
reg g1258;
reg g1259;
reg g1260;
reg g1251;
reg g1252;
reg g1253;
reg g1254;
reg g1176;
reg g1161;
reg g1168;
reg g1172;
reg g1173;
reg g1174;
reg g1175;
reg g1142;
reg g1145;
reg g1148;
reg g1164;
reg g1165;
reg g1166;
reg g1167;
reg g1171;
reg g1151;
reg g1152;
reg g1155;
reg g1158;
reg g1214;
reg g1221;
reg g1228;
reg g1229;
reg g1230;
reg g1234;
reg g1235;
reg g1186;
reg g1244;
reg g1245;
reg g1262;
reg g1263;
reg g1261;
reg g1265;
reg g1266;
reg g1264;
reg g1268;
reg g1269;
reg g1267;
reg g1271;
reg g1272;
reg g1270;
reg g1273;
reg g1276;
reg g1279;
reg g1282;
reg g1285;
reg g1288;
reg g1300;
reg g1303;
reg g1306;
reg g1291;
reg g1294;
reg g1297;
reg g1177;
reg g1180;
reg g1183;
reg g1192;
reg g1193;
reg g1194;
reg g1195;
reg g1200;
reg g1201;
reg g1202;
reg g1203;
reg g1204;
reg g1205;
reg g1206;
reg g1211;
reg g1215;
reg g1216;
reg g1217;
reg g1218;
reg g1219;
reg g1220;
reg g1222;
reg g1223;
reg g1224;
reg g1227;
reg g1309;
reg g1312;
reg g1315;
reg g1316;
reg g1345;
reg g1326;
reg g1319;
reg g1339;
reg g1332;
reg g1346;
reg g1358;
reg g1352;
reg g1365;
reg g1372;
reg g1378;
reg g1385;
reg g1386;
reg g1384;
reg g1388;
reg g1389;
reg g1387;
reg g1391;
reg g1392;
reg g1390;
reg g1394;
reg g1395;
reg g1393;
reg g1397;
reg g1398;
reg g1396;
reg g1400;
reg g1401;
reg g1399;
reg g1403;
reg g1404;
reg g1402;
reg g1406;
reg g1407;
reg g1405;
reg g1409;
reg g1410;
reg g1408;
reg g1412;
reg g1413;
reg g1411;
reg g1415;
reg g1416;
reg g1414;
reg g1418;
reg g1419;
reg g1417;
reg g1421;
reg g1422;
reg g1420;
reg g1424;
reg g1425;
reg g1423;
reg g1520;
reg g1517;
reg g1547;
reg g1512;
reg g1513;
reg g1511;
reg g1515;
reg g1516;
reg g1514;
reg g1524;
reg g1525;
reg g1523;
reg g1527;
reg g1528;
reg g1526;
reg g1530;
reg g1531;
reg g1529;
reg g1533;
reg g1534;
reg g1532;
reg g1536;
reg g1537;
reg g1535;
reg g1539;
reg g1540;
reg g1538;
reg g1542;
reg g1543;
reg g1541;
reg g1545;
reg g1546;
reg g1544;
reg g1551;
reg g1552;
reg g1550;
reg g1554;
reg g1555;
reg g1553;
reg g1557;
reg g1558;
reg g1556;
reg g1560;
reg g1561;
reg g1559;
reg g1567;
reg g1570;
reg g1573;
reg g1612;
reg g1615;
reg g1618;
reg g1576;
reg g1579;
reg g1582;
reg g1621;
reg g1624;
reg g1627;
reg g1585;
reg g1588;
reg g1591;
reg g1630;
reg g1633;
reg g1636;
reg g1594;
reg g1597;
reg g1600;
reg g1639;
reg g1642;
reg g1645;
reg g1603;
reg g1606;
reg g1609;
reg g1648;
reg g1651;
reg g1654;
reg g1466;
reg g1462;
reg g1457;
reg g1453;
reg g1448;
reg g1444;
reg g1439;
reg g1435;
reg g1430;
reg g1426;
reg g1562;
reg g1564;
reg g1563;
reg g1657;
reg g1786;
reg g1782;
reg g1690;
reg g1735;
reg g1724;
reg g1727;
reg g1750;
reg g1739;
reg g1742;
reg g1765;
reg g1754;
reg g1757;
reg g1779;
reg g1769;
reg g1772;
reg g1789;
reg g1792;
reg g1795;
reg g1798;
reg g1801;
reg g1804;
reg g1808;
reg g1809;
reg g1807;
reg g1810;
reg g1813;
reg g1816;
reg g1819;
reg g1822;
reg g1825;
reg g1829;
reg g1830;
reg g1828;
reg g1693;
reg g1694;
reg g1695;
reg g1696;
reg g1697;
reg g1698;
reg g1699;
reg g1700;
reg g1701;
reg g1703;
reg g1704;
reg g1702;
reg g1784;
reg g1785;
reg g1783;
reg g1831;
reg g1832;
reg g1833;
reg g1834;
reg g1835;
reg g1660;
reg g1661;
reg g1662;
reg g1663;
reg g1664;
reg g1665;
reg g1666;
reg g1667;
reg g1668;
reg g1669;
reg g1670;
reg g1671;
reg g1672;
reg g1680;
reg g1686;
reg g1689;
reg g1678;
reg g1677;
reg g1676;
reg g1675;
reg g1685;
reg g1684;
reg g1683;
reg g1682;
reg g1681;
reg g1679;
reg g1723;
reg g1730;
reg g1731;
reg g1732;
reg g1733;
reg g1734;
reg g1738;
reg g1745;
reg g1746;
reg g1747;
reg g1748;
reg g1749;
reg g1753;
reg g1760;
reg g1761;
reg g1762;
reg g1763;
reg g1764;
reg g1768;
reg g1775;
reg g1776;
reg g1777;
reg g1778;
reg g1705;
reg g1706;
reg g1712;
reg g1718;
reg g1925;
reg g1931;
reg g1930;
reg g1934;
reg g1937;
reg g1890;
reg g1893;
reg g1903;
reg g1904;
reg g1944;
reg g1949;
reg g1950;
reg g1951;
reg g1952;
reg g1953;
reg g1954;
reg g1945;
reg g1946;
reg g1947;
reg g1948;
reg g1870;
reg g1855;
reg g1862;
reg g1866;
reg g1867;
reg g1868;
reg g1869;
reg g1836;
reg g1839;
reg g1842;
reg g1858;
reg g1859;
reg g1860;
reg g1861;
reg g1865;
reg g1845;
reg g1846;
reg g1849;
reg g1852;
reg g1908;
reg g1915;
reg g1922;
reg g1923;
reg g1924;
reg g1928;
reg g1929;
reg g1880;
reg g1938;
reg g1939;
reg g1956;
reg g1957;
reg g1955;
reg g1959;
reg g1960;
reg g1958;
reg g1962;
reg g1963;
reg g1961;
reg g1965;
reg g1966;
reg g1964;
reg g1967;
reg g1970;
reg g1973;
reg g1976;
reg g1979;
reg g1982;
reg g1994;
reg g1997;
reg g2000;
reg g1985;
reg g1988;
reg g1991;
reg g1871;
reg g1874;
reg g1877;
reg g1886;
reg g1887;
reg g1888;
reg g1889;
reg g1894;
reg g1895;
reg g1896;
reg g1897;
reg g1898;
reg g1899;
reg g1900;
reg g1905;
reg g1909;
reg g1910;
reg g1911;
reg g1912;
reg g1913;
reg g1914;
reg g1916;
reg g1917;
reg g1918;
reg g1921;
reg g2003;
reg g2006;
reg g2009;
reg g2010;
reg g2039;
reg g2020;
reg g2013;
reg g2033;
reg g2026;
reg g2040;
reg g2052;
reg g2046;
reg g2059;
reg g2066;
reg g2072;
reg g2079;
reg g2080;
reg g2078;
reg g2082;
reg g2083;
reg g2081;
reg g2085;
reg g2086;
reg g2084;
reg g2088;
reg g2089;
reg g2087;
reg g2091;
reg g2092;
reg g2090;
reg g2094;
reg g2095;
reg g2093;
reg g2097;
reg g2098;
reg g2096;
reg g2100;
reg g2101;
reg g2099;
reg g2103;
reg g2104;
reg g2102;
reg g2106;
reg g2107;
reg g2105;
reg g2109;
reg g2110;
reg g2108;
reg g2112;
reg g2113;
reg g2111;
reg g2115;
reg g2116;
reg g2114;
reg g2118;
reg g2119;
reg g2117;
reg g2214;
reg g2211;
reg g2241;
reg g2206;
reg g2207;
reg g2205;
reg g2209;
reg g2210;
reg g2208;
reg g2218;
reg g2219;
reg g2217;
reg g2221;
reg g2222;
reg g2220;
reg g2224;
reg g2225;
reg g2223;
reg g2227;
reg g2228;
reg g2226;
reg g2230;
reg g2231;
reg g2229;
reg g2233;
reg g2234;
reg g2232;
reg g2236;
reg g2237;
reg g2235;
reg g2239;
reg g2240;
reg g2238;
reg g2245;
reg g2246;
reg g2244;
reg g2248;
reg g2249;
reg g2247;
reg g2251;
reg g2252;
reg g2250;
reg g2254;
reg g2255;
reg g2253;
reg g2261;
reg g2264;
reg g2267;
reg g2306;
reg g2309;
reg g2312;
reg g2270;
reg g2273;
reg g2276;
reg g2315;
reg g2318;
reg g2321;
reg g2279;
reg g2282;
reg g2285;
reg g2324;
reg g2327;
reg g2330;
reg g2288;
reg g2291;
reg g2294;
reg g2333;
reg g2336;
reg g2339;
reg g2297;
reg g2300;
reg g2303;
reg g2342;
reg g2345;
reg g2348;
reg g2160;
reg g2156;
reg g2151;
reg g2147;
reg g2142;
reg g2138;
reg g2133;
reg g2129;
reg g2124;
reg g2120;
reg g2256;
reg g2258;
reg g2257;
reg g2351;
reg g2480;
reg g2476;
reg g2384;
reg g2429;
reg g2418;
reg g2421;
reg g2444;
reg g2433;
reg g2436;
reg g2459;
reg g2448;
reg g2451;
reg g2473;
reg g2463;
reg g2466;
reg g2483;
reg g2486;
reg g2489;
reg g2492;
reg g2495;
reg g2498;
reg g2502;
reg g2503;
reg g2501;
reg g2504;
reg g2507;
reg g2510;
reg g2513;
reg g2516;
reg g2519;
reg g2523;
reg g2524;
reg g2522;
reg g2387;
reg g2388;
reg g2389;
reg g2390;
reg g2391;
reg g2392;
reg g2393;
reg g2394;
reg g2395;
reg g2397;
reg g2398;
reg g2396;
reg g2478;
reg g2479;
reg g2477;
reg g2525;
reg g2526;
reg g2527;
reg g2528;
reg g2529;
reg g2354;
reg g2355;
reg g2356;
reg g2357;
reg g2358;
reg g2359;
reg g2360;
reg g2361;
reg g2362;
reg g2363;
reg g2364;
reg g2365;
reg g2366;
reg g2374;
reg g2380;
reg g2383;
reg g2372;
reg g2371;
reg g2370;
reg g2369;
reg g2379;
reg g2378;
reg g2377;
reg g2376;
reg g2375;
reg g2373;
reg g2417;
reg g2424;
reg g2425;
reg g2426;
reg g2427;
reg g2428;
reg g2432;
reg g2439;
reg g2440;
reg g2441;
reg g2442;
reg g2443;
reg g2447;
reg g2454;
reg g2455;
reg g2456;
reg g2457;
reg g2458;
reg g2462;
reg g2469;
reg g2470;
reg g2471;
reg g2472;
reg g2399;
reg g2400;
reg g2406;
reg g2412;
reg g2619;
reg g2625;
reg g2624;
reg g2628;
reg g2631;
reg g2584;
reg g2587;
reg g2597;
reg g2598;
reg g2638;
reg g2643;
reg g2644;
reg g2645;
reg g2646;
reg g2647;
reg g2648;
reg g2639;
reg g2640;
reg g2641;
reg g2642;
reg g2564;
reg g2549;
reg g2556;
reg g2560;
reg g2561;
reg g2562;
reg g2563;
reg g2530;
reg g2533;
reg g2536;
reg g2552;
reg g2553;
reg g2554;
reg g2555;
reg g2559;
reg g2539;
reg g2540;
reg g2543;
reg g2546;
reg g2602;
reg g2609;
reg g2616;
reg g2617;
reg g2618;
reg g2622;
reg g2623;
reg g2574;
reg g2632;
reg g2633;
reg g2650;
reg g2651;
reg g2649;
reg g2653;
reg g2654;
reg g2652;
reg g2656;
reg g2657;
reg g2655;
reg g2659;
reg g2660;
reg g2658;
reg g2661;
reg g2664;
reg g2667;
reg g2670;
reg g2673;
reg g2676;
reg g2688;
reg g2691;
reg g2694;
reg g2679;
reg g2682;
reg g2685;
reg g2565;
reg g2568;
reg g2571;
reg g2580;
reg g2581;
reg g2582;
reg g2583;
reg g2588;
reg g2589;
reg g2590;
reg g2591;
reg g2592;
reg g2593;
reg g2594;
reg g2599;
reg g2603;
reg g2604;
reg g2605;
reg g2606;
reg g2607;
reg g2608;
reg g2610;
reg g2611;
reg g2612;
reg g2615;
reg g2697;
reg g2700;
reg g2703;
reg g2704;
reg g2733;
reg g2714;
reg g2707;
reg g2727;
reg g2720;
reg g2734;
reg g2746;
reg g2740;
reg g2753;
reg g2760;
reg g2766;
reg g2773;
reg g2774;
reg g2772;
reg g2776;
reg g2777;
reg g2775;
reg g2779;
reg g2780;
reg g2778;
reg g2782;
reg g2783;
reg g2781;
reg g2785;
reg g2786;
reg g2784;
reg g2788;
reg g2789;
reg g2787;
reg g2791;
reg g2792;
reg g2790;
reg g2794;
reg g2795;
reg g2793;
reg g2797;
reg g2798;
reg g2796;
reg g2800;
reg g2801;
reg g2799;
reg g2803;
reg g2804;
reg g2802;
reg g2806;
reg g2807;
reg g2805;
reg g2809;
reg g2810;
reg g2808;
reg g2812;
reg g2813;
reg g2811;
reg g3054;
reg g3079;
reg g3080;
reg g3043;
reg g3044;
reg g3045;
reg g3046;
reg g3047;
reg g3048;
reg g3049;
reg g3050;
reg g3051;
reg g3052;
reg g3053;
reg g3055;
reg g3056;
reg g3057;
reg g3058;
reg g3059;
reg g3060;
reg g3061;
reg g3062;
reg g3063;
reg g3064;
reg g3065;
reg g3066;
reg g3067;
reg g3068;
reg g3069;
reg g3070;
reg g3071;
reg g3072;
reg g3073;
reg g3074;
reg g3075;
reg g3076;
reg g3077;
reg g3078;
reg g2997;
reg g2993;
reg g2998;
reg g3006;
reg g3002;
reg g3013;
reg g3010;
reg g3024;
reg g3018;
reg g3028;
reg g3036;
reg g3032;
reg g3040;
reg g2986;
reg g2987;
reg g48;
reg g45;
reg g42;
reg g39;
reg g27;
reg g30;
reg g33;
reg g36;
reg g3083;
reg g26;
reg g2992;
reg g23;
reg g20;
reg g17;
reg g11;
reg g14;
reg g5;
reg g8;
reg g2;
reg g2990;
reg g2991;
reg g1;
wire g18281;
wire g20592;
wire g29827;
wire g16081;
wire g24124;
wire g17318;
wire g29394;
wire II30149;
wire g13447;
wire g30503;
wire g22225;
wire g24850;
wire II39056;
wire g23625;
wire II22919;
wire g10306;
wire g17674;
wire g13491;
wire g28911;
wire g14745;
wire g28845;
wire g30086;
wire g24831;
wire g24362;
wire g8508;
wire g6136;
wire II14712;
wire g30484;
wire g10300;
wire II14615;
wire II37128;
wire g11145;
wire g29928;
wire II30754;
wire g26774;
wire II20550;
wire g27059;
wire g26797;
wire g30797;
wire g20649;
wire g16015;
wire g26716;
wire g6426;
wire g10764;
wire g26734;
wire g8932;
wire II32535;
wire g22800;
wire II29448;
wire g13576;
wire g24396;
wire g19524;
wire g6045;
wire II25037;
wire II36234;
wire II18509;
wire g30716;
wire g24600;
wire g25379;
wire II32323;
wire g5845;
wire II28792;
wire II16965;
wire g22712;
wire g20454;
wire g3250;
wire g13626;
wire g22527;
wire II21908;
wire g28160;
wire g7600;
wire II35964;
wire II27335;
wire II21819;
wire g27547;
wire g24903;
wire g21458;
wire II40137;
wire g26632;
wire g17865;
wire g22719;
wire g21081;
wire g8862;
wire g4136;
wire g8938;
wire g5913;
wire g23609;
wire II29372;
wire g18644;
wire II29125;
wire g9034;
wire g25907;
wire II18100;
wire g22735;
wire II32851;
wire g23150;
wire g15647;
wire g28840;
wire g22695;
wire g7521;
wire g29308;
wire II25855;
wire g19900;
wire g10560;
wire g29740;
wire g24742;
wire g22314;
wire g21780;
wire g12193;
wire II22282;
wire g25200;
wire g22036;
wire g29098;
wire II34017;
wire II25857;
wire g19765;
wire II32695;
wire II18314;
wire g17694;
wire II21793;
wire II25820;
wire II33686;
wire II17200;
wire g22220;
wire g29295;
wire II34818;
wire g23556;
wire II29522;
wire g28186;
wire II36311;
wire II20514;
wire gbuf3;
wire g9635;
wire II22527;
wire g28168;
wire g10783;
wire g23276;
wire g28773;
wire g28619;
wire g29301;
wire g10230;
wire g19449;
wire g21375;
wire g17729;
wire II40101;
wire g23536;
wire g27065;
wire g14327;
wire II40832;
wire g21615;
wire g10495;
wire g27481;
wire g19638;
wire g10186;
wire II17730;
wire g30816;
wire g29873;
wire g22625;
wire g6015;
wire g20573;
wire II26642;
wire g15809;
wire g23984;
wire g4939;
wire II29656;
wire II18136;
wire g21135;
wire g18334;
wire II40209;
wire g8885;
wire g16039;
wire g21117;
wire g19028;
wire g14764;
wire g11650;
wire g22269;
wire g6101;
wire g23183;
wire g24906;
wire g20420;
wire g29336;
wire g30376;
wire g28925;
wire g30833;
wire g8123;
wire g4854;
wire g25630;
wire g9109;
wire g11565;
wire g16045;
wire g12868;
wire II15882;
wire II29145;
wire g4919;
wire g25413;
wire II38178;
wire II14489;
wire g30608;
wire g16066;
wire g8817;
wire II23667;
wire g11907;
wire II21674;
wire g18465;
wire II29399;
wire g23297;
wire g17652;
wire g11584;
wire g18048;
wire II23645;
wire g23313;
wire g13413;
wire g8704;
wire g13171;
wire g14158;
wire g22284;
wire g15520;
wire II36379;
wire II33596;
wire g21876;
wire g10270;
wire II17919;
wire II19794;
wire g6142;
wire II36993;
wire g30219;
wire II36690;
wire g28052;
wire g5989;
wire g19903;
wire II40706;
wire g29575;
wire g5363;
wire g12921;
wire g13642;
wire g20790;
wire g3931;
wire g5185;
wire g15179;
wire g27523;
wire g11900;
wire II20526;
wire II36601;
wire g29151;
wire g17136;
wire g10217;
wire g23051;
wire II21313;
wire g25232;
wire II29675;
wire g10117;
wire II20476;
wire g20273;
wire II23207;
wire g30946;
wire g19156;
wire g22142;
wire II34722;
wire g29246;
wire g28361;
wire g15593;
wire g16392;
wire g5935;
wire g27479;
wire g28059;
wire g15148;
wire II38339;
wire II35028;
wire g30646;
wire II35473;
wire g30764;
wire g22313;
wire g11811;
wire g20462;
wire g18994;
wire g14143;
wire g15989;
wire g20953;
wire II29694;
wire g30469;
wire g24796;
wire g21020;
wire g30333;
wire g12599;
wire II31769;
wire g26277;
wire g21550;
wire g30882;
wire g24519;
wire g18389;
wire g15210;
wire g30302;
wire g27138;
wire g10400;
wire II37665;
wire II37488;
wire II21249;
wire g26301;
wire II40288;
wire g22638;
wire g27184;
wire g8678;
wire II19542;
wire g20753;
wire g4699;
wire g12804;
wire g20496;
wire g10405;
wire g29957;
wire g22467;
wire g4168;
wire g28151;
wire g26806;
wire g4930;
wire II22924;
wire g4720;
wire g19314;
wire g12179;
wire II24539;
wire g24446;
wire g12485;
wire g24565;
wire II22845;
wire g29362;
wire g16881;
wire II39324;
wire g28344;
wire g30746;
wire II28494;
wire II31772;
wire g13194;
wire g21524;
wire g9582;
wire g10099;
wire g26480;
wire g24149;
wire g22246;
wire g25279;
wire g30491;
wire g13656;
wire g15720;
wire g7962;
wire g26606;
wire g19843;
wire g24069;
wire g5305;
wire II13962;
wire II33858;
wire II32453;
wire g17637;
wire g17252;
wire g26448;
wire g17704;
wire g14114;
wire g17090;
wire g13047;
wire II18232;
wire g15867;
wire g24427;
wire II17373;
wire g16345;
wire g16179;
wire II23894;
wire II40218;
wire g5971;
wire g11731;
wire g12041;
wire g11169;
wire g4702;
wire g13138;
wire g25781;
wire g8556;
wire g10201;
wire g29948;
wire g12122;
wire g4064;
wire g20836;
wire g26045;
wire g8250;
wire g19312;
wire g20789;
wire g16991;
wire g20614;
wire g10453;
wire II22900;
wire II35000;
wire g22117;
wire g30228;
wire II33278;
wire g18803;
wire II17992;
wire g18531;
wire g7856;
wire g8257;
wire g11344;
wire g30245;
wire II39541;
wire g24300;
wire g23917;
wire g17954;
wire g27575;
wire II33828;
wire g26357;
wire II34980;
wire g16767;
wire g16788;
wire g16446;
wire g11506;
wire g27693;
wire II26726;
wire g26667;
wire II16270;
wire g30689;
wire g10328;
wire g5815;
wire g25106;
wire II28169;
wire g29485;
wire g9289;
wire II26440;
wire g13477;
wire g27401;
wire II27228;
wire g17901;
wire g12217;
wire g22276;
wire g13366;
wire II20592;
wire II21563;
wire II30823;
wire g19668;
wire g27756;
wire g11045;
wire g7646;
wire g5210;
wire g30986;
wire g24003;
wire g26416;
wire g17143;
wire g18954;
wire II27119;
wire g19023;
wire g15602;
wire II16203;
wire II38459;
wire g25032;
wire g25946;
wire g24088;
wire g30265;
wire II29357;
wire g25131;
wire g5142;
wire g11759;
wire g8159;
wire g7896;
wire g29996;
wire g18286;
wire II24716;
wire g20342;
wire II18617;
wire II18461;
wire g10373;
wire II35425;
wire g8293;
wire g15304;
wire II36420;
wire g18917;
wire g11745;
wire g18003;
wire g14371;
wire g30550;
wire II13158;
wire g10969;
wire g23215;
wire g23563;
wire II19174;
wire II13775;
wire II19739;
wire II40200;
wire II13984;
wire g29973;
wire g16108;
wire g30682;
wire g30568;
wire g8915;
wire g3398;
wire II31496;
wire g24359;
wire g29257;
wire II22063;
wire g12233;
wire II38617;
wire g27904;
wire II29442;
wire II40484;
wire g10332;
wire II31670;
wire g30344;
wire g19142;
wire g27133;
wire g26145;
wire g30010;
wire II28594;
wire II16321;
wire g10007;
wire II32919;
wire II33633;
wire g30526;
wire g11550;
wire g24493;
wire g26614;
wire II26960;
wire g9111;
wire g7676;
wire II15256;
wire g30296;
wire g27508;
wire g18884;
wire g13559;
wire g24034;
wire g10854;
wire II22783;
wire g10333;
wire g26469;
wire g5894;
wire II25838;
wire g30403;
wire g26206;
wire II18211;
wire g13098;
wire g20133;
wire g30288;
wire g27422;
wire g10616;
wire g6029;
wire II40605;
wire II24292;
wire g12340;
wire g25977;
wire g28337;
wire g29175;
wire g27317;
wire g25627;
wire g29943;
wire II31784;
wire II25111;
wire g18656;
wire g24257;
wire g12505;
wire g19201;
wire II32159;
wire g5766;
wire g28211;
wire g22657;
wire II39157;
wire g4283;
wire g20526;
wire g23489;
wire g10165;
wire g30779;
wire II25606;
wire II34686;
wire II19412;
wire II18455;
wire g26872;
wire g16708;
wire II38807;
wire II23556;
wire g26826;
wire g14309;
wire g19861;
wire g11108;
wire g13373;
wire g8640;
wire g20307;
wire g14554;
wire g9919;
wire g25261;
wire g18811;
wire g25994;
wire g27298;
wire g30159;
wire g8844;
wire g27946;
wire g17157;
wire g13022;
wire g29288;
wire g18653;
wire g27794;
wire II19759;
wire gbuf130;
wire II35413;
wire g16733;
wire II24131;
wire g14060;
wire II31889;
wire g19192;
wire g11022;
wire II16062;
wire g29641;
wire g26697;
wire g23595;
wire g17248;
wire g6977;
wire g16074;
wire II18192;
wire g29340;
wire g25165;
wire g27590;
wire g21939;
wire g16484;
wire g26902;
wire g17219;
wire g29478;
wire g13219;
wire g13226;
wire g19282;
wire g13420;
wire g25596;
wire g24237;
wire g15251;
wire g22412;
wire g11324;
wire II15213;
wire gbuf35;
wire g21097;
wire g10729;
wire g27923;
wire II28019;
wire II15012;
wire g28220;
wire II19986;
wire II17889;
wire II32143;
wire II14195;
wire g19782;
wire g24846;
wire g21913;
wire II32189;
wire g27310;
wire g28612;
wire II18545;
wire II26377;
wire II27927;
wire g23863;
wire II13578;
wire g23476;
wire II40091;
wire g18188;
wire g23289;
wire g15562;
wire g13251;
wire g28761;
wire II37020;
wire II31056;
wire g19721;
wire gbuf211;
wire g10043;
wire g28524;
wire g10653;
wire g28903;
wire g23941;
wire II31802;
wire II17140;
wire g7709;
wire g7950;
wire II35856;
wire g28108;
wire g21211;
wire g27252;
wire g19720;
wire g8026;
wire g25833;
wire g23234;
wire II36486;
wire II27050;
wire g17597;
wire g20385;
wire II36250;
wire II37599;
wire g12005;
wire II40515;
wire g23974;
wire g17578;
wire g27772;
wire II37800;
wire g23433;
wire g22980;
wire II37965;
wire g29181;
wire g13428;
wire g17177;
wire g24973;
wire g12157;
wire II33813;
wire g29093;
wire g22196;
wire II25445;
wire g16265;
wire g7610;
wire g28177;
wire II32952;
wire g22750;
wire g19185;
wire II35548;
wire II34156;
wire g8490;
wire II24005;
wire g15118;
wire g9426;
wire II37011;
wire g20220;
wire II13239;
wire g19710;
wire g15747;
wire g29267;
wire g14059;
wire II36358;
wire II25089;
wire g25533;
wire II27014;
wire g24411;
wire II32892;
wire II41090;
wire g13498;
wire g26610;
wire II27008;
wire II24763;
wire g17212;
wire g21609;
wire II41114;
wire g19226;
wire g22045;
wire g23693;
wire g13540;
wire g15496;
wire g10463;
wire II38151;
wire II18731;
wire g23077;
wire g15997;
wire II18001;
wire g26572;
wire g9366;
wire g13610;
wire g12689;
wire II32074;
wire II19466;
wire g23410;
wire g8434;
wire II23966;
wire g18719;
wire g12775;
wire g12424;
wire g9048;
wire II38801;
wire II33482;
wire g18939;
wire g16351;
wire II19449;
wire II34830;
wire g23252;
wire g19289;
wire II23854;
wire II15629;
wire II34233;
wire g5829;
wire II35399;
wire g28804;
wire II16095;
wire g16426;
wire g19118;
wire II17837;
wire g25067;
wire g21476;
wire II31484;
wire gbuf121;
wire g15843;
wire II33504;
wire g21306;
wire g18726;
wire g27692;
wire II16918;
wire II39008;
wire g25057;
wire g8455;
wire g21032;
wire g15889;
wire g24014;
wire g28693;
wire g22204;
wire II17750;
wire g20516;
wire g21746;
wire II36705;
wire g29005;
wire II38737;
wire g30866;
wire gbuf23;
wire g22869;
wire g11876;
wire g28255;
wire g30521;
wire g22576;
wire g14703;
wire g19232;
wire g30677;
wire II21708;
wire g22147;
wire II34737;
wire g12847;
wire II21742;
wire g7869;
wire g20043;
wire g10102;
wire g11943;
wire g22179;
wire g29833;
wire II38951;
wire gbuf76;
wire g10175;
wire g19828;
wire g7358;
wire g7193;
wire g20311;
wire g30026;
wire g25667;
wire g30123;
wire g15603;
wire II25432;
wire g30593;
wire g20693;
wire g8531;
wire g26154;
wire g19982;
wire II36321;
wire g11222;
wire g19490;
wire II22581;
wire g15388;
wire II40600;
wire g15810;
wire g21751;
wire g19245;
wire g22606;
wire II25500;
wire g4094;
wire g26118;
wire g11884;
wire II36063;
wire g27086;
wire g11767;
wire II19404;
wire g27702;
wire g25967;
wire II29812;
wire g20895;
wire g13400;
wire g22186;
wire II34698;
wire g30382;
wire g26441;
wire g29638;
wire g27570;
wire g10880;
wire g15640;
wire II30026;
wire II18929;
wire g4611;
wire g11989;
wire g10918;
wire g29911;
wire g13432;
wire g22660;
wire g21226;
wire g20335;
wire g29515;
wire g10204;
wire g21268;
wire g11834;
wire g21970;
wire g17416;
wire II31115;
wire g8620;
wire g22948;
wire g18735;
wire g21812;
wire g12265;
wire II20909;
wire g4307;
wire g21823;
wire g11237;
wire II33611;
wire g23064;
wire g30061;
wire g24009;
wire II37291;
wire g12978;
wire g7926;
wire g15723;
wire g27907;
wire g24824;
wire g13853;
wire g26442;
wire g17630;
wire g23663;
wire g23459;
wire II26426;
wire g25758;
wire g24160;
wire g29661;
wire g15659;
wire g4395;
wire g11682;
wire II30350;
wire g19254;
wire g20053;
wire II40471;
wire g28242;
wire II40961;
wire g27119;
wire g21446;
wire g21846;
wire II26195;
wire g14573;
wire g30670;
wire g27435;
wire g6309;
wire g9758;
wire II14556;
wire g26753;
wire g10466;
wire g16479;
wire II23035;
wire g13075;
wire g18942;
wire g16091;
wire g3984;
wire II14631;
wire g4115;
wire g13356;
wire g25706;
wire II14574;
wire II40164;
wire g13816;
wire g23009;
wire g22458;
wire g23854;
wire g20406;
wire g10365;
wire g19971;
wire g28102;
wire g19803;
wire II33182;
wire g22549;
wire II22316;
wire g17556;
wire g5149;
wire g7538;
wire II37188;
wire g28472;
wire g5888;
wire g13518;
wire g20292;
wire II40254;
wire g17122;
wire g19808;
wire II39401;
wire g17042;
wire g25451;
wire II17054;
wire g28466;
wire II19952;
wire II18444;
wire g23627;
wire II24587;
wire g26835;
wire g15240;
wire II25580;
wire II23478;
wire g22154;
wire g15410;
wire g18850;
wire g26957;
wire II37885;
wire II23075;
wire II37459;
wire II22917;
wire II26574;
wire g19883;
wire g5326;
wire II18181;
wire II13232;
wire g30229;
wire g30963;
wire g24078;
wire g29761;
wire g25405;
wire g28997;
wire II38119;
wire g26882;
wire g11887;
wire II16303;
wire g9630;
wire g26240;
wire II25311;
wire II37379;
wire g25110;
wire g6066;
wire g18183;
wire g28381;
wire g26821;
wire g21335;
wire g30756;
wire g9936;
wire II28000;
wire g30949;
wire g25022;
wire g22705;
wire II32430;
wire g29464;
wire II30374;
wire II16653;
wire II38821;
wire g17878;
wire g10911;
wire II18677;
wire g16061;
wire II25655;
wire g12645;
wire g21040;
wire g5412;
wire g4409;
wire II30741;
wire g14882;
wire g29510;
wire g13280;
wire II22810;
wire g12328;
wire II20637;
wire g16863;
wire II40098;
wire g9766;
wire II28712;
wire g9160;
wire g24337;
wire II36411;
wire g21298;
wire g25019;
wire g11672;
wire g5400;
wire g17998;
wire g27236;
wire g10586;
wire II27232;
wire g25239;
wire g19597;
wire g20974;
wire g17012;
wire II22599;
wire g10599;
wire g10475;
wire g12197;
wire g4237;
wire g23052;
wire II29077;
wire g20157;
wire II37334;
wire g15494;
wire II38232;
wire g25655;
wire g15557;
wire g9257;
wire g23174;
wire g24180;
wire g26390;
wire II24205;
wire II13173;
wire g19932;
wire g23452;
wire II38725;
wire gbuf55;
wire g24098;
wire II14149;
wire g13805;
wire g27697;
wire II25733;
wire g22834;
wire g12172;
wire II19025;
wire g29431;
wire g12819;
wire II38958;
wire II37578;
wire g22810;
wire II35821;
wire g15827;
wire g13621;
wire II14538;
wire II23501;
wire g10935;
wire II35554;
wire g9442;
wire II38447;
wire II40784;
wire g26562;
wire II30598;
wire II19303;
wire g19042;
wire g29226;
wire g27315;
wire g17529;
wire g3238;
wire g24536;
wire g22451;
wire II40227;
wire II20532;
wire g30937;
wire g27747;
wire II38536;
wire g8341;
wire g27032;
wire g21354;
wire g10515;
wire g25253;
wire g14230;
wire g23746;
wire g10649;
wire g27466;
wire g11669;
wire II16930;
wire g21330;
wire II28249;
wire II23908;
wire g23579;
wire g22533;
wire g26686;
wire g26367;
wire II23191;
wire g29192;
wire II29016;
wire II36571;
wire g10255;
wire g5907;
wire g5835;
wire II18402;
wire g24588;
wire II16726;
wire g29508;
wire g19206;
wire g7906;
wire II15167;
wire g26022;
wire g10396;
wire g28316;
wire II24474;
wire g12024;
wire II35410;
wire II37137;
wire II21680;
wire g17021;
wire g27834;
wire g30371;
wire g29220;
wire g23512;
wire g11515;
wire g22676;
wire g15516;
wire g28249;
wire II17294;
wire g20098;
wire II14647;
wire g15873;
wire g16453;
wire g11051;
wire g24572;
wire II32422;
wire g22685;
wire II16309;
wire II21952;
wire g26083;
wire g10321;
wire g30854;
wire g11651;
wire g16986;
wire g26768;
wire II34400;
wire g15688;
wire g17018;
wire g22915;
wire II17895;
wire II30002;
wire g10679;
wire II16190;
wire g19736;
wire g17755;
wire g13297;
wire g8354;
wire II40475;
wire g13482;
wire g26428;
wire g24083;
wire g26006;
wire g27279;
wire II30908;
wire g29639;
wire g11188;
wire g27251;
wire II32492;
wire g13469;
wire g20333;
wire II23368;
wire g29436;
wire g17017;
wire g26062;
wire g28738;
wire g21083;
wire g22385;
wire II25672;
wire II18575;
wire g29781;
wire g17282;
wire g25151;
wire g15990;
wire II18082;
wire II41105;
wire II29291;
wire g29049;
wire g8690;
wire g19018;
wire g28141;
wire g19542;
wire II31724;
wire g21859;
wire g6421;
wire g28421;
wire g17682;
wire g10630;
wire g24037;
wire g30968;
wire g25770;
wire II32660;
wire g30828;
wire g21356;
wire g28439;
wire II13186;
wire g23245;
wire gbuf124;
wire g13969;
wire g16672;
wire II25597;
wire g13738;
wire g29556;
wire g24267;
wire g4948;
wire g19369;
wire II40107;
wire g7053;
wire g22092;
wire g27408;
wire g19351;
wire II35109;
wire g12376;
wire gbuf92;
wire II31426;
wire g23867;
wire g19648;
wire g19175;
wire g26640;
wire g12442;
wire g28078;
wire g20779;
wire g10512;
wire g10675;
wire II29478;
wire g28359;
wire g19874;
wire g18936;
wire II19784;
wire II35407;
wire g28834;
wire g16439;
wire g10294;
wire g15178;
wire g17161;
wire g29628;
wire g9100;
wire g3616;
wire g4035;
wire g29791;
wire g12078;
wire g5804;
wire II24678;
wire g5787;
wire g10639;
wire g21639;
wire g9894;
wire II33539;
wire g19699;
wire g27913;
wire g13134;
wire II15549;
wire g22885;
wire g20996;
wire II16185;
wire g27582;
wire g26282;
wire g19704;
wire g19972;
wire II15359;
wire g28007;
wire II16785;
wire g23310;
wire II24554;
wire g24243;
wire g22588;
wire II31841;
wire g30019;
wire g27002;
wire g28552;
wire g4662;
wire II37228;
wire g29283;
wire g11707;
wire g12108;
wire g28859;
wire g11762;
wire II37973;
wire g28069;
wire g18898;
wire II31562;
wire g5170;
wire g27271;
wire g10825;
wire g16829;
wire g26450;
wire g19560;
wire g15546;
wire g14234;
wire g19476;
wire g11069;
wire II38342;
wire II33532;
wire g9873;
wire g13243;
wire g25933;
wire g21819;
wire g8577;
wire g24897;
wire g8065;
wire g19884;
wire II23791;
wire g6227;
wire g24310;
wire g30030;
wire gbuf43;
wire II29610;
wire g21946;
wire II23880;
wire g19096;
wire II13228;
wire g8526;
wire II32704;
wire g13065;
wire g25983;
wire II33689;
wire g25827;
wire g20436;
wire g19277;
wire g9925;
wire II27328;
wire g10870;
wire g25419;
wire g5763;
wire II22667;
wire II35497;
wire II40110;
wire II21982;
wire g5041;
wire g24581;
wire g11059;
wire II31133;
wire II19891;
wire g8877;
wire g25699;
wire g10018;
wire g27228;
wire g15363;
wire g13368;
wire g10415;
wire g6000;
wire g20366;
wire g29703;
wire II24560;
wire g4564;
wire g25010;
wire II34111;
wire gbuf193;
wire II40724;
wire II21429;
wire g19270;
wire g26958;
wire II18488;
wire g25086;
wire g11216;
wire g13123;
wire II16172;
wire g7423;
wire g29270;
wire g12904;
wire g10036;
wire g21180;
wire g30724;
wire g27973;
wire II18527;
wire g9228;
wire g13033;
wire g28656;
wire II37716;
wire g22645;
wire II21609;
wire g13835;
wire g11785;
wire g13701;
wire g10147;
wire g28281;
wire II38278;
wire g20425;
wire g22875;
wire g9722;
wire g24938;
wire g10378;
wire g27729;
wire g6099;
wire g18788;
wire II15779;
wire g8382;
wire g11537;
wire g30392;
wire II19855;
wire g24859;
wire g24378;
wire g29736;
wire g28123;
wire g9355;
wire II24308;
wire g22754;
wire g16008;
wire g18649;
wire g19851;
wire g9027;
wire g17258;
wire II21329;
wire II40245;
wire g24386;
wire II31205;
wire g21599;
wire II27565;
wire g28678;
wire g20920;
wire II38920;
wire g28349;
wire g27820;
wire g26708;
wire g12932;
wire g20185;
wire g7795;
wire g11573;
wire g11501;
wire g30058;
wire g19238;
wire II38088;
wire g24208;
wire g15711;
wire g26815;
wire g28581;
wire g12531;
wire g24371;
wire II16472;
wire g29965;
wire g13052;
wire g26869;
wire g15757;
wire g29143;
wire g30361;
wire g23301;
wire g25289;
wire g26566;
wire g22650;
wire g8018;
wire g5982;
wire g8944;
wire g24782;
wire II33498;
wire II35058;
wire g8909;
wire II38172;
wire g24841;
wire II34579;
wire II35373;
wire g20901;
wire g14895;
wire g12691;
wire g29936;
wire g24223;
wire g17486;
wire g20644;
wire II18740;
wire II35035;
wire g5552;
wire g27414;
wire g18991;
wire II24500;
wire g16198;
wire g26609;
wire g26173;
wire g21012;
wire II38668;
wire II31937;
wire g11956;
wire g22363;
wire II37729;
wire II24123;
wire g21106;
wire g5949;
wire g14794;
wire II20586;
wire g13460;
wire II28201;
wire g5668;
wire g7528;
wire II35003;
wire g25147;
wire g14298;
wire II36598;
wire II36499;
wire g25123;
wire g8856;
wire g23182;
wire g13486;
wire g24475;
wire II30011;
wire II33399;
wire g15354;
wire II15836;
wire II40919;
wire g26019;
wire g12708;
wire II27146;
wire g6230;
wire II30161;
wire g29347;
wire g25124;
wire g25215;
wire g12186;
wire g29421;
wire g27540;
wire g24778;
wire g27288;
wire g16494;
wire g10269;
wire g17050;
wire g22841;
wire g29563;
wire g10260;
wire g17785;
wire g22774;
wire g15635;
wire g25388;
wire II18799;
wire g25029;
wire g17531;
wire g29685;
wire g21234;
wire g25688;
wire g23129;
wire g21362;
wire II27942;
wire II35083;
wire g21074;
wire g27200;
wire g10470;
wire g17148;
wire g15718;
wire g10661;
wire g26477;
wire II15833;
wire g8197;
wire g5706;
wire g24431;
wire II39164;
wire II40715;
wire g28923;
wire g22192;
wire g24053;
wire II29435;
wire g24406;
wire II23760;
wire II29007;
wire g10258;
wire g8485;
wire II37659;
wire g7576;
wire g26232;
wire g20780;
wire g10319;
wire g8467;
wire II40916;
wire g30974;
wire g27455;
wire II14413;
wire II27358;
wire g7878;
wire g19045;
wire g27207;
wire g26658;
wire g7549;
wire g20455;
wire g20345;
wire II40651;
wire g21903;
wire g16359;
wire g28661;
wire g11864;
wire g13127;
wire g14222;
wire g20285;
wire g16024;
wire g28192;
wire g21122;
wire II29142;
wire II26916;
wire II20848;
wire II37946;
wire g23408;
wire II26383;
wire g25664;
wire g13026;
wire g28073;
wire g10754;
wire g17351;
wire g11736;
wire II14478;
wire g19759;
wire g29316;
wire g27661;
wire g30478;
wire g5227;
wire II37296;
wire g24367;
wire II33402;
wire g21850;
wire g19795;
wire g25681;
wire g27071;
wire II23152;
wire II22981;
wire g30326;
wire g19940;
wire g8488;
wire II19852;
wire II20562;
wire g12438;
wire g18368;
wire g5776;
wire g26165;
wire g28237;
wire II37814;
wire II25880;
wire g14182;
wire g15263;
wire g26726;
wire II36516;
wire g24763;
wire g10949;
wire g9623;
wire g28025;
wire g16358;
wire g6032;
wire II29301;
wire g15890;
wire g28477;
wire g8141;
wire II33646;
wire II18206;
wire g27303;
wire g15174;
wire g26037;
wire g15296;
wire II40212;
wire g11199;
wire g4549;
wire II25234;
wire g27196;
wire g12876;
wire II38205;
wire g21965;
wire II35727;
wire g10813;
wire II29533;
wire g17717;
wire g10154;
wire II38524;
wire II31745;
wire g26120;
wire g30105;
wire II28119;
wire g9903;
wire g26644;
wire g16460;
wire g27266;
wire g26239;
wire II29317;
wire g16389;
wire g10316;
wire g12815;
wire g24921;
wire II31282;
wire g25227;
wire g23170;
wire g8518;
wire g27937;
wire g24522;
wire II37113;
wire II21809;
wire g27281;
wire g22077;
wire II40955;
wire g27683;
wire g28110;
wire g28680;
wire g27802;
wire g25589;
wire g30460;
wire II24992;
wire g14863;
wire g28413;
wire g26158;
wire g9174;
wire II25489;
wire g21870;
wire g26855;
wire gbuf164;
wire g21261;
wire g5675;
wire g5058;
wire g11796;
wire II23144;
wire g27105;
wire g18909;
wire gbuf188;
wire g11256;
wire II30359;
wire g27419;
wire g21665;
wire g12112;
wire g26860;
wire g24342;
wire II32686;
wire II39936;
wire g14957;
wire g20927;
wire g11190;
wire II30769;
wire II18019;
wire g13303;
wire g11998;
wire II36755;
wire II32847;
wire g15314;
wire g11933;
wire g25053;
wire g18968;
wire g25194;
wire g29118;
wire g11297;
wire II24696;
wire II35334;
wire g21618;
wire II25355;
wire g27345;
wire g10843;
wire g29771;
wire g5012;
wire g28839;
wire g8563;
wire II25782;
wire g5256;
wire g27980;
wire g25738;
wire g29565;
wire g6189;
wire g21894;
wire g30563;
wire g27075;
wire g23068;
wire g30887;
wire g10792;
wire II36630;
wire g25062;
wire g27535;
wire g24182;
wire II37740;
wire g22727;
wire g28687;
wire g30525;
wire g25075;
wire g4406;
wire g17737;
wire g21222;
wire g14205;
wire g8400;
wire g13204;
wire g16188;
wire II15915;
wire g25072;
wire g8212;
wire g21411;
wire II30748;
wire g13148;
wire g22796;
wire g18458;
wire g30119;
wire g21152;
wire II27488;
wire g5407;
wire II23172;
wire g28498;
wire g13346;
wire g14752;
wire II26796;
wire g12852;
wire g29776;
wire g19978;
wire II41065;
wire g16546;
wire g10106;
wire II21304;
wire II39368;
wire g28259;
wire g28607;
wire g11411;
wire g24804;
wire g20968;
wire g5745;
wire g12051;
wire g20433;
wire II19240;
wire II30362;
wire g17850;
wire g17150;
wire II25890;
wire g29756;
wire g23049;
wire g20919;
wire g13273;
wire II32583;
wire g29666;
wire g27024;
wire II30813;
wire g8631;
wire g9038;
wire g11800;
wire g21490;
wire g27706;
wire g19191;
wire g24147;
wire g24444;
wire g17128;
wire g20539;
wire g14776;
wire g12506;
wire g28212;
wire g21983;
wire g11971;
wire g29704;
wire g9062;
wire g29164;
wire g22143;
wire II38591;
wire g25796;
wire II39625;
wire g20084;
wire II29459;
wire g17223;
wire g18827;
wire g24413;
wire II34716;
wire g30253;
wire II29582;
wire g26783;
wire II17645;
wire g24233;
wire g19623;
wire II35737;
wire g30890;
wire II24325;
wire g12611;
wire g22183;
wire g16382;
wire g18897;
wire g21497;
wire II38330;
wire g5880;
wire g23610;
wire g14011;
wire g20586;
wire II34827;
wire g7841;
wire g29426;
wire g16583;
wire g19912;
wire g8276;
wire II30047;
wire g18415;
wire g13001;
wire g27604;
wire g11855;
wire g15578;
wire II30386;
wire g11599;
wire g22250;
wire g4845;
wire g11979;
wire g29353;
wire g9199;
wire g27504;
wire g9920;
wire II22715;
wire g13456;
wire g23524;
wire g10061;
wire g9081;
wire II19648;
wire g13503;
wire II35488;
wire g26222;
wire gbuf84;
wire II16071;
wire II16068;
wire g10525;
wire II30143;
wire g11048;
wire g26814;
wire II39361;
wire II38059;
wire II23218;
wire g30899;
wire g28982;
wire g8924;
wire II28727;
wire g30810;
wire II39815;
wire g19592;
wire II23911;
wire g23012;
wire g15701;
wire g30512;
wire g24276;
wire II16031;
wire g28199;
wire g14378;
wire II31640;
wire g7916;
wire II32595;
wire g25158;
wire g21219;
wire II34785;
wire g22546;
wire g21491;
wire g13864;
wire II39270;
wire g13290;
wire g7140;
wire g20379;
wire II33511;
wire g27595;
wire g30004;
wire II38211;
wire II34803;
wire g19390;
wire II31667;
wire II32365;
wire II25412;
wire g18578;
wire II16499;
wire g9450;
wire g15065;
wire g7141;
wire g27246;
wire II26874;
wire g15880;
wire g8997;
wire g27191;
wire II17311;
wire II34405;
wire g26790;
wire g22445;
wire II28470;
wire g12533;
wire II13113;
wire g26691;
wire II35141;
wire g11008;
wire g26055;
wire II23256;
wire II40799;
wire II26895;
wire g23770;
wire g14975;
wire g22559;
wire II18091;
wire g7661;
wire g22591;
wire g29807;
wire g11543;
wire g28434;
wire g23911;
wire II22657;
wire II30704;
wire g30915;
wire g13111;
wire g7877;
wire g6084;
wire II18199;
wire II25195;
wire g29234;
wire g23738;
wire II25406;
wire g19562;
wire II19510;
wire II40054;
wire II18114;
wire g21321;
wire g16804;
wire g11611;
wire g25360;
wire g10386;
wire g22512;
wire II27416;
wire g11827;
wire II30632;
wire g12346;
wire II16796;
wire g20392;
wire g25510;
wire II36147;
wire II33445;
wire g21343;
wire g30897;
wire II22705;
wire g21056;
wire II30173;
wire II20062;
wire g28935;
wire II17771;
wire g26316;
wire g23074;
wire g5260;
wire g16309;
wire g22176;
wire g18906;
wire g12324;
wire II37152;
wire II31574;
wire II31529;
wire g20625;
wire g17511;
wire g30337;
wire II36591;
wire g19326;
wire g29130;
wire g22065;
wire g24305;
wire g3248;
wire g11695;
wire g10592;
wire g17749;
wire g28099;
wire g28230;
wire g18290;
wire II18695;
wire II39333;
wire g19617;
wire g24112;
wire g20477;
wire g5822;
wire II30654;
wire g23570;
wire g22560;
wire g16846;
wire g11361;
wire g30448;
wire g7591;
wire g30823;
wire g20117;
wire g16472;
wire II39121;
wire g12752;
wire g28023;
wire g25339;
wire II30395;
wire g30859;
wire g30279;
wire II27402;
wire g16323;
wire g26068;
wire g14884;
wire g25183;
wire II37167;
wire g11453;
wire II23421;
wire g7809;
wire g9765;
wire g19674;
wire g27143;
wire II35817;
wire g12998;
wire g25383;
wire g5757;
wire II25985;
wire g5375;
wire g22739;
wire g21805;
wire g15506;
wire g30008;
wire g25036;
wire g24812;
wire g10626;
wire g7079;
wire II36954;
wire II26990;
wire g24179;
wire II20791;
wire II15955;
wire g10746;
wire g22123;
wire g22934;
wire II39859;
wire II36779;
wire g6184;
wire II30077;
wire g19384;
wire g24165;
wire g16619;
wire II33864;
wire g8559;
wire g27687;
wire g13324;
wire g26264;
wire II27900;
wire g17969;
wire g18975;
wire II19523;
wire g19079;
wire g4228;
wire g27256;
wire g30956;
wire g19695;
wire II30869;
wire g5279;
wire II27143;
wire g27558;
wire g19758;
wire g8542;
wire g22635;
wire g19381;
wire g22364;
wire g29045;
wire g30249;
wire g16230;
wire g30262;
wire g20619;
wire g29544;
wire g25332;
wire II28093;
wire g18523;
wire g22764;
wire g12282;
wire g26457;
wire g19155;
wire g8074;
wire g7769;
wire g12419;
wire g10808;
wire g10079;
wire g30544;
wire g11916;
wire g21640;
wire II40629;
wire g29496;
wire g22131;
wire g13564;
wire II16276;
wire g4354;
wire g23196;
wire g25135;
wire g24356;
wire g26107;
wire g30269;
wire g22236;
wire g28720;
wire g19196;
wire g21076;
wire g21881;
wire g30924;
wire g24451;
wire g10558;
wire g8666;
wire gbuf50;
wire g18837;
wire g12970;
wire g22294;
wire g30651;
wire g22558;
wire g30584;
wire g8983;
wire g18838;
wire II18187;
wire g13714;
wire II29960;
wire II18130;
wire g4379;
wire g26854;
wire g12385;
wire g21006;
wire II31706;
wire g6190;
wire g26538;
wire g20602;
wire II22989;
wire g20673;
wire II14822;
wire gbuf118;
wire g25000;
wire g19014;
wire g22105;
wire g13737;
wire g5714;
wire II34662;
wire g23791;
wire II20802;
wire g26213;
wire II21554;
wire II36438;
wire g18923;
wire g5422;
wire g5991;
wire g22002;
wire g25366;
wire g16252;
wire g13187;
wire g8102;
wire II24207;
wire g15467;
wire g18868;
wire II29619;
wire g12306;
wire g29282;
wire g30733;
wire II35783;
wire II23904;
wire g27498;
wire g22353;
wire g27214;
wire g15033;
wire g21889;
wire g16736;
wire g26620;
wire g12518;
wire g29458;
wire g16513;
wire g8448;
wire g19178;
wire g24833;
wire g12915;
wire g15786;
wire II25711;
wire II24351;
wire g28716;
wire II40191;
wire g27516;
wire g19070;
wire II13820;
wire II30586;
wire g25249;
wire II18055;
wire II22518;
wire II15354;
wire II16532;
wire g9883;
wire II26505;
wire g13381;
wire II37474;
wire g13154;
wire g24951;
wire II29632;
wire g17336;
wire II40444;
wire II31171;
wire II38518;
wire g25349;
wire gbuf185;
wire g28695;
wire II36882;
wire g22379;
wire g25856;
wire II40931;
wire II37757;
wire g24542;
wire g19924;
wire g24681;
wire g10123;
wire g22828;
wire II16338;
wire g20011;
wire II41099;
wire g26383;
wire g16725;
wire g18141;
wire g27099;
wire g13989;
wire g24218;
wire g28954;
wire II36909;
wire g16694;
wire g9121;
wire g7949;
wire g24091;
wire g27115;
wire g20322;
wire II33984;
wire g30801;
wire g24920;
wire g11662;
wire g27124;
wire II30738;
wire g27090;
wire gbuf74;
wire g28500;
wire g25311;
wire g22785;
wire g11351;
wire II30962;
wire g23330;
wire II22676;
wire g18406;
wire g30358;
wire g12463;
wire II24339;
wire II40083;
wire II13131;
wire g15847;
wire g20556;
wire g26985;
wire II16296;
wire g28267;
wire g26944;
wire g20522;
wire g24219;
wire g12990;
wire g17942;
wire II30233;
wire II32391;
wire g30223;
wire g24456;
wire gbuf157;
wire g10192;
wire II18332;
wire g19088;
wire g4433;
wire g15320;
wire g21488;
wire g26478;
wire g19032;
wire g24852;
wire g5417;
wire g29137;
wire II25078;
wire II16056;
wire g13851;
wire g30087;
wire g18983;
wire II36314;
wire g25814;
wire g22611;
wire g12476;
wire g8097;
wire g23022;
wire g20998;
wire g18218;
wire II25061;
wire g14767;
wire g28068;
wire g7779;
wire II33364;
wire II27200;
wire g25363;
wire g21312;
wire g24753;
wire g21214;
wire g25463;
wire II33016;
wire II24253;
wire g3365;
wire II26282;
wire g19778;
wire II17429;
wire II15890;
wire II14571;
wire g4959;
wire g11559;
wire II34916;
wire g19769;
wire g11213;
wire II27158;
wire g26866;
wire g8996;
wire g17082;
wire g8549;
wire II37197;
wire g22732;
wire g30933;
wire II18866;
wire g26406;
wire g9793;
wire g23197;
wire II25897;
wire g17582;
wire g26997;
wire g15920;
wire g28298;
wire g14614;
wire II37647;
wire g7802;
wire g23115;
wire g11842;
wire II14009;
wire g19111;
wire g28301;
wire g21453;
wire g7974;
wire II24613;
wire g24093;
wire II36915;
wire g13797;
wire g22970;
wire g17085;
wire g30691;
wire g13935;
wire g21647;
wire gbuf173;
wire g27715;
wire g23593;
wire g13687;
wire g23033;
wire g12456;
wire g8430;
wire g21007;
wire g26970;
wire g30029;
wire g22309;
wire g19345;
wire g4740;
wire g11899;
wire g5856;
wire g12312;
wire II17081;
wire g8575;
wire g19329;
wire II38245;
wire g24546;
wire II16225;
wire g17616;
wire g27007;
wire g8478;
wire g19555;
wire II25308;
wire gbuf119;
wire g20620;
wire g10839;
wire II25762;
wire g18115;
wire II20441;
wire g25808;
wire g15852;
wire g10924;
wire g20278;
wire g8443;
wire g18152;
wire g25282;
wire g17058;
wire g26308;
wire g30480;
wire g11702;
wire g21046;
wire g5621;
wire g30876;
wire II23999;
wire II37203;
wire g29402;
wire g15785;
wire II13098;
wire II40587;
wire g27269;
wire g20911;
wire g26761;
wire II35841;
wire g23684;
wire g29291;
wire g29528;
wire g30342;
wire II15616;
wire g13443;
wire gbuf33;
wire II14378;
wire g21164;
wire g13061;
wire g20136;
wire g21175;
wire g24862;
wire g19661;
wire g12099;
wire II24601;
wire g18270;
wire g24596;
wire II13149;
wire II25344;
wire II29513;
wire gbuf198;
wire g27839;
wire g27850;
wire II23639;
wire II40985;
wire g29918;
wire II24481;
wire g27018;
wire g11721;
wire g25209;
wire g16995;
wire g4058;
wire g21501;
wire II30254;
wire g24777;
wire g15830;
wire II16101;
wire gbuf17;
wire g23089;
wire II32509;
wire g8784;
wire II24150;
wire g12833;
wire II17486;
wire g23429;
wire g10725;
wire II22759;
wire II30639;
wire g15396;
wire g5849;
wire g13118;
wire g11776;
wire g30364;
wire g29538;
wire g29072;
wire g12759;
wire II40973;
wire II30791;
wire II37994;
wire g27046;
wire II29209;
wire II40886;
wire II23266;
wire g24691;
wire g16458;
wire g29924;
wire II24745;
wire g10583;
wire II18686;
wire g9133;
wire II30194;
wire g16282;
wire g25342;
wire g26800;
wire g4515;
wire II24317;
wire g17114;
wire g19602;
wire g29522;
wire g25599;
wire g11890;
wire II28065;
wire II15794;
wire g20610;
wire II18076;
wire g9774;
wire g23587;
wire g12481;
wire g29206;
wire g16017;
wire g26202;
wire g17301;
wire II25320;
wire g11287;
wire g24315;
wire g27154;
wire g12440;
wire g4970;
wire g20658;
wire g12412;
wire g7826;
wire II40664;
wire g28640;
wire II34012;
wire II28148;
wire g12146;
wire g29581;
wire g5390;
wire II36441;
wire g16131;
wire g10183;
wire g20567;
wire g29266;
wire g11370;
wire II40435;
wire g19125;
wire g18928;
wire II17737;
wire g27360;
wire g22987;
wire II33909;
wire g23602;
wire g8613;
wire II39539;
wire g17993;
wire g17710;
wire g19678;
wire II25495;
wire g12101;
wire g13550;
wire II13904;
wire g25950;
wire g27052;
wire g20063;
wire g11692;
wire g30930;
wire g22715;
wire II24368;
wire II21577;
wire g25143;
wire II36781;
wire g23715;
wire g21731;
wire g18089;
wire g12245;
wire g5084;
wire g23205;
wire g30804;
wire g4480;
wire g18708;
wire g9676;
wire g26003;
wire II14882;
wire g17758;
wire II19862;
wire g16289;
wire g23768;
wire g19816;
wire g16138;
wire g7999;
wire g9893;
wire g16134;
wire II28876;
wire g4685;
wire II17849;
wire g22945;
wire g13525;
wire g22033;
wire g28555;
wire g30783;
wire g28336;
wire g11995;
wire g10498;
wire g25990;
wire II18683;
wire g28705;
wire g26683;
wire g29502;
wire g8176;
wire II24280;
wire II14544;
wire g15897;
wire II17846;
wire II38028;
wire g29654;
wire II22884;
wire g23679;
wire II38632;
wire g29818;
wire g24463;
wire II25004;
wire g11386;
wire g7724;
wire II30272;
wire II33831;
wire g23264;
wire g10451;
wire II32443;
wire g11629;
wire II33737;
wire g12292;
wire g15664;
wire II33882;
wire g29388;
wire g7329;
wire II29249;
wire g11965;
wire II34118;
wire g29724;
wire g8755;
wire g12223;
wire g28350;
wire g26364;
wire g28746;
wire g8570;
wire II24452;
wire g11873;
wire g22165;
wire g10522;
wire II33561;
wire g18224;
wire g23845;
wire II27110;
wire II36948;
wire g13740;
wire g25157;
wire II27243;
wire g15480;
wire g30658;
wire II34026;
wire II14049;
wire g28080;
wire II35777;
wire II21256;
wire II28210;
wire II25682;
wire g28701;
wire II30519;
wire g28273;
wire g10012;
wire II27182;
wire g27323;
wire g8395;
wire g8719;
wire g5975;
wire g5397;
wire g26961;
wire II39347;
wire g29120;
wire II29484;
wire g3960;
wire g28897;
wire g19571;
wire g16749;
wire g24106;
wire g28485;
wire g25978;
wire g21775;
wire g26592;
wire g17165;
wire g8161;
wire g20357;
wire g16050;
wire II38606;
wire g13952;
wire II17936;
wire II18969;
wire II18163;
wire g20946;
wire g20937;
wire II18737;
wire g25745;
wire g17949;
wire II21822;
wire g12353;
wire g28081;
wire g7785;
wire g18755;
wire g29415;
wire g27235;
wire g21035;
wire g18120;
wire g9090;
wire II17925;
wire II13849;
wire g22939;
wire g7685;
wire g12054;
wire II34433;
wire g5912;
wire g12952;
wire g7389;
wire g18876;
wire g30836;
wire II24387;
wire g23377;
wire g28036;
wire II36942;
wire g6713;
wire II14496;
wire g9302;
wire g25140;
wire II31868;
wire g29696;
wire g15851;
wire g19665;
wire II21340;
wire gbuf65;
wire II40787;
wire g13332;
wire g30775;
wire g3338;
wire g28305;
wire II36404;
wire g27571;
wire II19195;
wire g18552;
wire g23161;
wire II37961;
wire g22272;
wire g8350;
wire g5605;
wire g16104;
wire g8659;
wire g20389;
wire II31931;
wire g24176;
wire II15429;
wire II40167;
wire g18912;
wire II23163;
wire g10457;
wire II22718;
wire II40441;
wire g21605;
wire II31853;
wire II34755;
wire g30120;
wire g29133;
wire g24328;
wire g11928;
wire II30868;
wire g22949;
wire g23112;
wire g29008;
wire g3995;
wire g27467;
wire g15691;
wire g20904;
wire g29784;
wire g12213;
wire g30109;
wire g19146;
wire g7560;
wire g21244;
wire g25274;
wire g13495;
wire g4289;
wire II37775;
wire g12524;
wire g16908;
wire gbuf26;
wire g29660;
wire g10251;
wire g21339;
wire g19730;
wire g18958;
wire II28365;
wire g23214;
wire g13139;
wire g10519;
wire II29194;
wire g8421;
wire II33529;
wire II36156;
wire g21157;
wire II23504;
wire g18950;
wire g12994;
wire g29313;
wire g24441;
wire g12782;
wire g29952;
wire II18004;
wire II26497;
wire g28734;
wire g4304;
wire g18469;
wire II36693;
wire g24623;
wire g13175;
wire II27149;
wire g15133;
wire g19749;
wire II36933;
wire g16183;
wire II24363;
wire II20820;
wire g29571;
wire g27295;
wire g25401;
wire II15912;
wire II25099;
wire II40997;
wire II18572;
wire g30982;
wire g17215;
wire g14291;
wire g23272;
wire g5890;
wire g13011;
wire g27028;
wire g8636;
wire g30649;
wire g18880;
wire g18652;
wire II25243;
wire g30407;
wire g23485;
wire g10642;
wire g29550;
wire II30032;
wire g30283;
wire g10003;
wire II39909;
wire g30187;
wire II21626;
wire g22555;
wire II16684;
wire II32178;
wire II34779;
wire g26693;
wire g19654;
wire g20718;
wire g5224;
wire g6170;
wire II26695;
wire II37796;
wire II21165;
wire g11802;
wire g8859;
wire g11883;
wire g6116;
wire II40032;
wire g24286;
wire g10101;
wire g11385;
wire II25666;
wire II39469;
wire g28970;
wire g27314;
wire g23105;
wire g29148;
wire g19846;
wire g24612;
wire g25265;
wire g15048;
wire g11347;
wire g12004;
wire g24253;
wire g10850;
wire g23970;
wire g18648;
wire II37394;
wire II25351;
wire g4263;
wire II25126;
wire II23860;
wire II40524;
wire II38386;
wire g17715;
wire g26840;
wire g26553;
wire g20227;
wire II36283;
wire II14027;
wire g4912;
wire g24898;
wire II22786;
wire g28065;
wire g8022;
wire g27927;
wire g24144;
wire g24365;
wire g24842;
wire II36711;
wire g18206;
wire g7540;
wire g30442;
wire g17797;
wire g26374;
wire II30215;
wire g19726;
wire g30132;
wire g26619;
wire g26209;
wire II24464;
wire g4538;
wire g24559;
wire g4809;
wire g4979;
wire g4788;
wire g5263;
wire g17221;
wire g18435;
wire II16630;
wire g5241;
wire g3460;
wire g11278;
wire g5825;
wire II40122;
wire g28098;
wire g24388;
wire g24605;
wire g12289;
wire g24497;
wire II27399;
wire g28137;
wire g25216;
wire g13423;
wire II17363;
wire g26731;
wire g29253;
wire g29305;
wire g12252;
wire II16117;
wire g4592;
wire g22041;
wire g26877;
wire g19451;
wire II38421;
wire g16370;
wire g9115;
wire II31493;
wire II37629;
wire g28171;
wire g23871;
wire g19007;
wire g16488;
wire g24552;
wire g28979;
wire g10056;
wire g4250;
wire g14130;
wire g29082;
wire II38683;
wire g22503;
wire II35545;
wire g20429;
wire g15638;
wire g29260;
wire g20269;
wire g27527;
wire II29500;
wire g27021;
wire II23695;
wire g9782;
wire g8336;
wire g15672;
wire g23284;
wire II16166;
wire II19996;
wire II40805;
wire II26664;
wire g9407;
wire g26576;
wire g9519;
wire II32982;
wire g22744;
wire II29168;
wire II16247;
wire g26260;
wire g20732;
wire g17173;
wire g28990;
wire II33520;
wire g23413;
wire II13110;
wire g23826;
wire g18679;
wire II26231;
wire g17439;
wire g25949;
wire g11265;
wire g18441;
wire g29992;
wire g20766;
wire g26178;
wire g23238;
wire g24747;
wire II24966;
wire g22851;
wire g21390;
wire II15623;
wire II32156;
wire g13389;
wire II18370;
wire II30041;
wire g28224;
wire II38148;
wire II32409;
wire II38710;
wire g23945;
wire g21113;
wire g13163;
wire g22336;
wire II37260;
wire II40307;
wire II40925;
wire g29709;
wire g23567;
wire II20794;
wire g5107;
wire g12369;
wire II25325;
wire g28652;
wire g26832;
wire g10980;
wire g24478;
wire g20088;
wire g4447;
wire II36407;
wire II13221;
wire g4038;
wire g6019;
wire gbuf200;
wire II25198;
wire g20942;
wire g10169;
wire g19222;
wire g23135;
wire II16759;
wire II31799;
wire g4766;
wire II35319;
wire g14459;
wire II32548;
wire g9725;
wire II13275;
wire g28966;
wire II37901;
wire g8852;
wire g21489;
wire g3978;
wire g18744;
wire g13190;
wire II33879;
wire II39124;
wire g22200;
wire g30322;
wire g5917;
wire g30022;
wire II32922;
wire g9127;
wire g13053;
wire g11830;
wire g4339;
wire II39376;
wire II33870;
wire g30812;
wire g17856;
wire g15631;
wire g30488;
wire g26702;
wire g27779;
wire g11727;
wire g30055;
wire g5952;
wire II27137;
wire g19647;
wire g26712;
wire g15017;
wire g10886;
wire II32081;
wire g22262;
wire g10932;
wire II39385;
wire II38122;
wire gbuf150;
wire II13990;
wire g19753;
wire II36582;
wire g20542;
wire g22300;
wire g20470;
wire g10397;
wire II13215;
wire II32561;
wire g17734;
wire g10219;
wire g24902;
wire g27751;
wire g28844;
wire g5416;
wire g5306;
wire g21064;
wire g17342;
wire II40490;
wire g8514;
wire g24513;
wire g24561;
wire g28778;
wire II35297;
wire g24392;
wire g27454;
wire g28412;
wire II36423;
wire II37356;
wire g19681;
wire II34680;
wire II18317;
wire g21227;
wire g22266;
wire II37608;
wire g13537;
wire II22875;
wire g27427;
wire g25082;
wire II18335;
wire g13435;
wire II34353;
wire II20601;
wire g25128;
wire II19482;
wire g12843;
wire II33807;
wire II36585;
wire II38007;
wire g17048;
wire gbuf190;
wire II18506;
wire II18417;
wire g23473;
wire g10096;
wire g10676;
wire g27748;
wire g29624;
wire gbuf114;
wire g27705;
wire II14900;
wire II31298;
wire g26679;
wire g27562;
wire g5677;
wire II20649;
wire II16018;
wire II14113;
wire II25429;
wire g8284;
wire g13905;
wire g16033;
wire g15274;
wire g16836;
wire g12808;
wire g22360;
wire g14390;
wire g15323;
wire g28480;
wire g5378;
wire g5182;
wire g5731;
wire g11813;
wire II32335;
wire g22310;
wire g18519;
wire g10087;
wire g21099;
wire II22813;
wire g10021;
wire g28164;
wire g9065;
wire II31244;
wire g22998;
wire g28041;
wire II30134;
wire g19628;
wire g13404;
wire g20981;
wire II40462;
wire II21415;
wire g29823;
wire g13093;
wire g24909;
wire II15800;
wire g24993;
wire g21566;
wire g26345;
wire II22640;
wire II39770;
wire g19943;
wire II13943;
wire g27181;
wire II14624;
wire g25942;
wire II21720;
wire II32913;
wire II24475;
wire g29117;
wire II34689;
wire g24525;
wire II13320;
wire g18843;
wire g17724;
wire g9613;
wire g6832;
wire II13119;
wire II32526;
wire g13397;
wire g28393;
wire g26738;
wire g19552;
wire g22691;
wire II39466;
wire g19718;
wire g6031;
wire g28406;
wire g19848;
wire g21102;
wire g5772;
wire g29958;
wire g28055;
wire II34071;
wire g27567;
wire g18352;
wire g22288;
wire II29030;
wire g19318;
wire g25228;
wire II40275;
wire g26587;
wire g11904;
wire II16200;
wire II28184;
wire g17465;
wire g29357;
wire g25119;
wire g24533;
wire g5818;
wire II15526;
wire g15577;
wire g30713;
wire g27475;
wire g5286;
wire g4671;
wire II40257;
wire g28377;
wire II18392;
wire g19605;
wire g27485;
wire g29249;
wire g10401;
wire II27041;
wire g10225;
wire g17464;
wire g20576;
wire g28117;
wire g13071;
wire g10540;
wire II38199;
wire g26041;
wire g15144;
wire g19152;
wire g20487;
wire g19058;
wire g30334;
wire g26819;
wire g16070;
wire g7009;
wire g30704;
wire II26416;
wire II37252;
wire g11028;
wire g17670;
wire g3878;
wire II35849;
wire II33545;
wire g5719;
wire g24281;
wire g23394;
wire g23292;
wire g15403;
wire g21142;
wire II18016;
wire g8329;
wire g28367;
wire g8708;
wire II24677;
wire g10080;
wire II13999;
wire II39791;
wire g27737;
wire g27150;
wire II31130;
wire g28877;
wire g25231;
wire g13233;
wire g29397;
wire g29327;
wire g5954;
wire II27733;
wire II18250;
wire g11496;
wire g19761;
wire g8934;
wire II37614;
wire g13340;
wire g29242;
wire g13942;
wire II18692;
wire g21181;
wire g9911;
wire g14486;
wire g10210;
wire g22281;
wire g13339;
wire g7581;
wire g26558;
wire g19952;
wire g8866;
wire g29332;
wire g23553;
wire II25174;
wire g19907;
wire II16697;
wire g30096;
wire g29577;
wire g27083;
wire g5145;
wire g5811;
wire II17027;
wire g10865;
wire g28294;
wire g8560;
wire II26528;
wire g16841;
wire g22582;
wire g6145;
wire g27061;
wire II14897;
wire g21554;
wire g18699;
wire g11809;
wire g10078;
wire g30849;
wire g21793;
wire II20500;
wire g8014;
wire g28348;
wire g23155;
wire g12321;
wire g8254;
wire g4861;
wire g16445;
wire g22517;
wire II33469;
wire g5163;
wire g26765;
wire g28826;
wire g23999;
wire g23776;
wire g18453;
wire II23715;
wire g30743;
wire g20247;
wire II17203;
wire II21813;
wire g5934;
wire g10325;
wire g29932;
wire g18337;
wire g21863;
wire g19748;
wire g12083;
wire g11734;
wire g27733;
wire g19559;
wire g26639;
wire g21452;
wire g11741;
wire g19211;
wire g14115;
wire II38752;
wire II40116;
wire g21720;
wire g30537;
wire g23265;
wire g6025;
wire g18997;
wire g30479;
wire g20416;
wire g8832;
wire g15175;
wire II39325;
wire gbuf161;
wire g28145;
wire g8150;
wire g29370;
wire g18346;
wire g29687;
wire g4174;
wire II25117;
wire g22701;
wire g8552;
wire II24522;
wire g26079;
wire g28936;
wire g10433;
wire II37787;
wire g27900;
wire g13913;
wire II15553;
wire g10818;
wire g16018;
wire g29552;
wire g12561;
wire g26465;
wire g26087;
wire g25031;
wire g30341;
wire g19181;
wire II22671;
wire g19637;
wire g10392;
wire g16298;
wire II36462;
wire g29815;
wire II33006;
wire II38740;
wire g26594;
wire II18476;
wire g13625;
wire g20094;
wire II13169;
wire g26423;
wire II32479;
wire g19731;
wire II18429;
wire II32410;
wire g16386;
wire g17100;
wire g20599;
wire g28467;
wire g17779;
wire g7697;
wire g10075;
wire II25691;
wire g14724;
wire g10015;
wire g26743;
wire g30495;
wire II27897;
wire g10628;
wire g4298;
wire II30191;
wire g23335;
wire g25749;
wire II29238;
wire g8635;
wire g28228;
wire g23582;
wire g21736;
wire g8828;
wire II19865;
wire g30858;
wire g24584;
wire g12789;
wire II32708;
wire g17451;
wire g5121;
wire g21779;
wire II18139;
wire g9427;
wire g27167;
wire g24027;
wire II31490;
wire g27679;
wire g14630;
wire g19195;
wire g10682;
wire II30269;
wire g6425;
wire g8180;
wire g25717;
wire g25132;
wire g30579;
wire II39933;
wire g23716;
wire g21353;
wire g14006;
wire II24372;
wire g10645;
wire II13680;
wire II25159;
wire g21447;
wire g28855;
wire g16632;
wire g17523;
wire II23235;
wire g21010;
wire g14525;
wire g15160;
wire g26796;
wire g12104;
wire g21049;
wire II28488;
wire g30268;
wire II19576;
wire g5592;
wire g26080;
wire g28178;
wire g5832;
wire g15442;
wire g30668;
wire II29013;
wire g21580;
wire g19479;
wire g30901;
wire II14917;
wire II36513;
wire g24323;
wire g23042;
wire g24125;
wire g29923;
wire II21852;
wire g17046;
wire II39982;
wire II30689;
wire II16538;
wire g24407;
wire II23460;
wire II21772;
wire g22396;
wire II28582;
wire g23742;
wire g16089;
wire g14558;
wire g28425;
wire g28215;
wire gbuf95;
wire g27838;
wire g27188;
wire g16953;
wire g30908;
wire II24291;
wire g15034;
wire II40572;
wire g13104;
wire g4746;
wire g13089;
wire g20562;
wire II15276;
wire g27372;
wire gbuf136;
wire g28358;
wire II21420;
wire g29691;
wire g24261;
wire g27990;
wire g29795;
wire g5735;
wire g19530;
wire g19061;
wire II28755;
wire g28285;
wire g30083;
wire g11120;
wire g30452;
wire II30941;
wire g10710;
wire g15475;
wire g29171;
wire g27012;
wire g12446;
wire g11766;
wire II34815;
wire II24752;
wire g12908;
wire II32696;
wire g22804;
wire g18988;
wire II34761;
wire g15814;
wire II17928;
wire g27147;
wire g22381;
wire gbuf128;
wire g25354;
wire II39895;
wire g28900;
wire g29081;
wire g19001;
wire g8873;
wire g28312;
wire II19872;
wire g6188;
wire g23249;
wire g13298;
wire g10290;
wire II17786;
wire g14001;
wire II24632;
wire g30052;
wire g28727;
wire g15246;
wire g7353;
wire g8794;
wire g13042;
wire II21787;
wire II14499;
wire II34728;
wire II15345;
wire g27449;
wire g5398;
wire g24989;
wire g29915;
wire g5427;
wire II34710;
wire g6058;
wire g11867;
wire II18220;
wire II32940;
wire g21636;
wire II18689;
wire g4476;
wire g9105;
wire g14212;
wire II37575;
wire g30674;
wire g9957;
wire II15308;
wire g29390;
wire g13705;
wire II22881;
wire g29369;
wire II32609;
wire g30014;
wire g22328;
wire II33652;
wire g7346;
wire g19015;
wire g27586;
wire g13069;
wire g25015;
wire II35491;
wire g14342;
wire II38220;
wire g23849;
wire g20368;
wire II35686;
wire g10424;
wire g27855;
wire g10207;
wire II16176;
wire g11055;
wire II40478;
wire g16290;
wire g4516;
wire II31778;
wire g30374;
wire g8745;
wire g21094;
wire II19932;
wire g12551;
wire g18902;
wire g29216;
wire g16571;
wire II35803;
wire g24304;
wire g5027;
wire g28364;
wire g30729;
wire g12222;
wire g28280;
wire g25240;
wire II40185;
wire g19128;
wire g5808;
wire g24881;
wire II16559;
wire g23624;
wire II16169;
wire g30387;
wire II22663;
wire II35530;
wire II31757;
wire g8810;
wire II40850;
wire g30179;
wire g7927;
wire g16011;
wire II34428;
wire g13347;
wire II30988;
wire g26578;
wire g12020;
wire g27328;
wire g8521;
wire g19097;
wire g16536;
wire II17206;
wire g25647;
wire g19785;
wire g8809;
wire g12494;
wire g13264;
wire g28455;
wire g20992;
wire g26327;
wire II19591;
wire g5800;
wire II36093;
wire g27342;
wire g20950;
wire II36786;
wire II30508;
wire g16042;
wire g11781;
wire g28355;
wire II21548;
wire II27209;
wire g13172;
wire g21427;
wire II31417;
wire g9390;
wire g29970;
wire II32994;
wire g13893;
wire II32997;
wire II29093;
wire II38038;
wire II16714;
wire II35673;
wire g30720;
wire II40152;
wire II17753;
wire II36752;
wire II24582;
wire g18629;
wire g25762;
wire g14228;
wire g16835;
wire g24357;
wire g8305;
wire g5683;
wire II37149;
wire II22998;
wire g26968;
wire g15339;
wire g4348;
wire II14644;
wire II21381;
wire g6041;
wire II32092;
wire g16417;
wire II18320;
wire g5323;
wire II38437;
wire g26244;
wire g21029;
wire II21479;
wire g10855;
wire II34180;
wire g29129;
wire II20414;
wire II27194;
wire g27799;
wire II14928;
wire g26346;
wire g24033;
wire g26980;
wire g10441;
wire II15593;
wire g24893;
wire g6637;
wire g16528;
wire gbuf180;
wire g28730;
wire g20450;
wire g4070;
wire g24234;
wire II29326;
wire g19249;
wire II28323;
wire g29473;
wire g10822;
wire g12478;
wire g23893;
wire g8535;
wire g20978;
wire g20697;
wire g21646;
wire II14945;
wire II15511;
wire g12271;
wire II38674;
wire g10367;
wire g24756;
wire g24700;
wire II20390;
wire g24950;
wire g15823;
wire g9886;
wire g6051;
wire II35136;
wire g13157;
wire g8827;
wire g24489;
wire g14098;
wire II15185;
wire II37017;
wire g19987;
wire g13229;
wire g22641;
wire II17834;
wire g28739;
wire g26445;
wire g26393;
wire g11603;
wire g26770;
wire g20682;
wire g7349;
wire g23059;
wire g25046;
wire g17634;
wire g9075;
wire II14868;
wire gbuf176;
wire II33304;
wire g21678;
wire II25801;
wire g10170;
wire II33961;
wire g17542;
wire II24445;
wire g26777;
wire g26215;
wire g27121;
wire II28009;
wire g23178;
wire g16243;
wire g28944;
wire II40643;
wire g21000;
wire g14520;
wire g8980;
wire g23835;
wire g25041;
wire g4383;
wire II20619;
wire II16110;
wire g27696;
wire g27265;
wire II19886;
wire II35933;
wire g20648;
wire g19250;
wire g10280;
wire g29110;
wire II24594;
wire g18430;
wire g19806;
wire g15655;
wire g18961;
wire g10910;
wire g16934;
wire II18827;
wire g7776;
wire II36749;
wire g19255;
wire g19820;
wire g28886;
wire g27559;
wire g21974;
wire g29155;
wire II29921;
wire g16423;
wire II18638;
wire g20439;
wire II30023;
wire g20057;
wire g13857;
wire g16965;
wire II38822;
wire II40772;
wire g30013;
wire II40988;
wire II19733;
wire g28299;
wire g25393;
wire gbuf79;
wire II15326;
wire g12460;
wire g30127;
wire g23165;
wire g25937;
wire g11428;
wire g16420;
wire g22621;
wire g21843;
wire II18854;
wire II19533;
wire g30352;
wire g12198;
wire II25848;
wire g12269;
wire g17345;
wire II18845;
wire g28251;
wire II37297;
wire g5221;
wire II23338;
wire g4614;
wire g14099;
wire II34321;
wire II27155;
wire II36224;
wire gbuf145;
wire g20093;
wire g24245;
wire II29369;
wire II26171;
wire g19335;
wire II19569;
wire g20690;
wire g26601;
wire g18727;
wire g10906;
wire g21254;
wire II38282;
wire gbuf51;
wire II25477;
wire g30215;
wire II40420;
wire g19541;
wire g21807;
wire g28064;
wire II40568;
wire g19051;
wire g27865;
wire g24577;
wire g10362;
wire g29138;
wire II27176;
wire g20885;
wire II23559;
wire II34165;
wire g11719;
wire g9749;
wire g26472;
wire g24529;
wire g16867;
wire II40811;
wire II18817;
wire g30635;
wire II25213;
wire g4555;
wire g25235;
wire g20025;
wire g22108;
wire II33507;
wire II30014;
wire g28015;
wire II32251;
wire II29525;
wire g16154;
wire g19951;
wire II18716;
wire II25228;
wire gbuf8;
wire g13398;
wire g28324;
wire II36612;
wire II29395;
wire II27278;
wire gbuf207;
wire II40634;
wire II32725;
wire g5970;
wire g24772;
wire g18313;
wire g28106;
wire g25988;
wire II24188;
wire g9773;
wire II36099;
wire g15198;
wire g20282;
wire g29518;
wire g12898;
wire g18169;
wire g5900;
wire II26913;
wire g28156;
wire g22216;
wire g19107;
wire g21402;
wire gbuf27;
wire II13959;
wire II24417;
wire g20876;
wire g18854;
wire g18998;
wire g13201;
wire II27920;
wire g10379;
wire g13220;
wire g30541;
wire g30082;
wire g6945;
wire g29765;
wire g25409;
wire g30752;
wire II30857;
wire g29489;
wire II25645;
wire II23219;
wire g19827;
wire g29468;
wire gbuf20;
wire II13801;
wire II34734;
wire II19833;
wire g30642;
wire g22599;
wire g18947;
wire g5355;
wire g13409;
wire g22153;
wire g20153;
wire gbuf42;
wire II33382;
wire g27484;
wire g27035;
wire g13252;
wire g5150;
wire g22830;
wire g11502;
wire g15794;
wire II21806;
wire g5008;
wire g16858;
wire g27843;
wire g12090;
wire II16258;
wire g19944;
wire g13234;
wire II19829;
wire g18603;
wire g22682;
wire g29744;
wire II23982;
wire g10596;
wire g21865;
wire g9150;
wire II26639;
wire II19777;
wire II15866;
wire g29057;
wire II29496;
wire g24480;
wire g17824;
wire II36897;
wire g19091;
wire g30594;
wire g23850;
wire g11315;
wire g26886;
wire g28374;
wire II17768;
wire g5005;
wire g29168;
wire g15856;
wire g27784;
wire II25050;
wire II31598;
wire g12452;
wire II24648;
wire g30481;
wire g19566;
wire g29616;
wire g22104;
wire g22083;
wire g21156;
wire g4437;
wire g16431;
wire g4688;
wire II34207;
wire g21271;
wire g20005;
wire g25071;
wire g22048;
wire g27349;
wire g17874;
wire g11647;
wire II23926;
wire g26352;
wire g24781;
wire g8029;
wire g6632;
wire g20002;
wire g19030;
wire g18096;
wire g27922;
wire g13391;
wire g13261;
wire g30436;
wire II40432;
wire g16647;
wire g13214;
wire II30278;
wire g11822;
wire II39945;
wire g19457;
wire g29032;
wire g22673;
wire g29186;
wire g9453;
wire g7638;
wire g29968;
wire II35975;
wire II24567;
wire g29276;
wire II17975;
wire II38866;
wire g10568;
wire g25095;
wire g20965;
wire g21399;
wire g6630;
wire II25867;
wire g29861;
wire g25305;
wire g20164;
wire g20819;
wire g5403;
wire g21302;
wire g29075;
wire II29019;
wire g11511;
wire II15262;
wire g13208;
wire g5944;
wire g12259;
wire g6080;
wire g26905;
wire II38462;
wire g25573;
wire II27017;
wire g22615;
wire g25198;
wire g13225;
wire g15800;
wire g23547;
wire g5749;
wire II28959;
wire g23611;
wire g20020;
wire g12499;
wire II21301;
wire II38620;
wire II40874;
wire g29422;
wire II32668;
wire g18987;
wire g8791;
wire g21890;
wire g23368;
wire g13144;
wire g7643;
wire g20371;
wire g27806;
wire II15902;
wire g27896;
wire g21172;
wire II23874;
wire II22687;
wire II36668;
wire g22793;
wire g21193;
wire II39761;
wire II15853;
wire II16814;
wire g10312;
wire g5884;
wire g29774;
wire g25370;
wire g28684;
wire g27987;
wire II26237;
wire g10157;
wire g6087;
wire g5423;
wire II38412;
wire g27555;
wire g26363;
wire g27255;
wire g12536;
wire g22114;
wire g16969;
wire g16718;
wire g20396;
wire g20964;
wire II20595;
wire g19483;
wire II36144;
wire II34656;
wire II24538;
wire g26792;
wire II36459;
wire g8964;
wire II31535;
wire g17265;
wire g20659;
wire g16523;
wire g16099;
wire g6036;
wire g19103;
wire g11666;
wire g29669;
wire g12161;
wire g23268;
wire g22171;
wire g18823;
wire g10284;
wire g21991;
wire II29912;
wire II25671;
wire g28430;
wire II22860;
wire II31457;
wire g24672;
wire g26248;
wire g23822;
wire g29344;
wire II17989;
wire g29717;
wire g29286;
wire g24877;
wire II14219;
wire g28492;
wire g24657;
wire II13937;
wire g30508;
wire g18308;
wire g16551;
wire II21137;
wire gbuf141;
wire g30102;
wire g30955;
wire g15791;
wire g7673;
wire g26007;
wire II35443;
wire g29237;
wire g27608;
wire II33415;
wire g27239;
wire g21410;
wire g24047;
wire g22422;
wire g13489;
wire g28132;
wire II29135;
wire g13860;
wire g19870;
wire II20589;
wire g15222;
wire II32904;
wire II27053;
wire II19415;
wire g20376;
wire g7688;
wire g11520;
wire g22254;
wire g17965;
wire II40796;
wire g25193;
wire g17249;
wire II32967;
wire g22654;
wire g15900;
wire g29646;
wire II16511;
wire II28189;
wire g20132;
wire g7594;
wire g21623;
wire g8928;
wire II17042;
wire g5252;
wire g14690;
wire g4023;
wire g17447;
wire II29978;
wire g28764;
wire II35416;
wire g16879;
wire II16123;
wire g27177;
wire g19235;
wire g30663;
wire g19879;
wire g10531;
wire g24272;
wire g28428;
wire II28743;
wire g28556;
wire II17765;
wire g22509;
wire II37155;
wire g17764;
wire g12894;
wire g25881;
wire g20113;
wire g25929;
wire g15741;
wire g18635;
wire g16054;
wire g15978;
wire g29230;
wire g13149;
wire II32469;
wire g24808;
wire g29449;
wire g16781;
wire g21249;
wire g5869;
wire g8906;
wire g18849;
wire g6367;
wire II37131;
wire g10772;
wire g21051;
wire g5587;
wire II41011;
wire g18478;
wire g20469;
wire II20839;
wire II32400;
wire II22604;
wire g19304;
wire II23277;
wire g25974;
wire gbuf131;
wire g21764;
wire g28390;
wire g28300;
wire g25623;
wire g28389;
wire g23636;
wire g29203;
wire II33583;
wire g20139;
wire g27241;
wire II21865;
wire II31121;
wire g27471;
wire g19242;
wire g24963;
wire g22168;
wire g25211;
wire II15992;
wire II23047;
wire g26670;
wire g11004;
wire II29559;
wire g30400;
wire g8752;
wire g25450;
wire II40994;
wire g30275;
wire g17079;
wire g13328;
wire g9924;
wire g22258;
wire g23574;
wire II19667;
wire g25997;
wire g26466;
wire II31188;
wire II36873;
wire g10892;
wire II16504;
wire II38226;
wire g18784;
wire g11556;
wire g17396;
wire g21369;
wire II23056;
wire g20362;
wire g18012;
wire II21461;
wire g12607;
wire II38832;
wire g22871;
wire II40016;
wire g29442;
wire g7476;
wire II15995;
wire g4389;
wire II14357;
wire g5369;
wire gbuf81;
wire II20486;
wire g14910;
wire g4735;
wire II35992;
wire g24070;
wire II19803;
wire g29069;
wire II38869;
wire g19356;
wire II40194;
wire g9003;
wire g10382;
wire g27531;
wire g17698;
wire g5615;
wire g21626;
wire II28509;
wire II14446;
wire g28494;
wire II31883;
wire g29620;
wire g7736;
wire II40934;
wire g26547;
wire g7479;
wire g12837;
wire g11699;
wire g8614;
wire g3244;
wire g24151;
wire II23403;
wire g11141;
wire g4791;
wire g21367;
wire g25684;
wire g21291;
wire II22797;
wire g9293;
wire g17144;
wire g16004;
wire g12115;
wire II24029;
wire g26397;
wire II17933;
wire g7799;
wire g30443;
wire g22068;
wire g9242;
wire g5877;
wire g19574;
wire g3306;
wire g16490;
wire II41018;
wire g27985;
wire g29961;
wire g21238;
wire g21502;
wire II16041;
wire g22866;
wire II38924;
wire g25323;
wire II16569;
wire g30862;
wire II35716;
wire g29681;
wire g14483;
wire g25223;
wire g22651;
wire II20033;
wire II26455;
wire g30258;
wire g19799;
wire g10538;
wire g9631;
wire g16992;
wire II35031;
wire g22358;
wire g11936;
wire II36627;
wire g11568;
wire g15837;
wire g30397;
wire g22128;
wire g29339;
wire g5962;
wire g23518;
wire g13654;
wire g30575;
wire g28277;
wire g5790;
wire II39130;
wire II25971;
wire g21070;
wire g22211;
wire g23299;
wire II35698;
wire g21160;
wire g13199;
wire g13046;
wire g22845;
wire g23000;
wire g5963;
wire g12943;
wire g28022;
wire II27593;
wire II33843;
wire II29288;
wire g29219;
wire g22583;
wire g30112;
wire g17773;
wire II35455;
wire II17807;
wire g22221;
wire II17860;
wire g23386;
wire II32576;
wire g21324;
wire g30793;
wire II37815;
wire g18893;
wire g15879;
wire g15714;
wire g17482;
wire g21611;
wire g26781;
wire II35756;
wire g7530;
wire g26313;
wire g26236;
wire II17951;
wire g5730;
wire g8386;
wire II24427;
wire g14119;
wire g8120;
wire g12194;
wire g27480;
wire g23803;
wire g22494;
wire g12153;
wire II24575;
wire gbuf103;
wire g30556;
wire g27842;
wire g21935;
wire II36066;
wire II24149;
wire g17476;
wire II30486;
wire g5862;
wire g25127;
wire II15239;
wire g15903;
wire II40534;
wire g24402;
wire g13257;
wire g21251;
wire II38428;
wire gbuf115;
wire g12553;
wire II30392;
wire g23907;
wire II38848;
wire g26648;
wire g17372;
wire g10672;
wire II37508;
wire g19789;
wire g23143;
wire II29122;
wire g30438;
wire g27101;
wire g25520;
wire g5795;
wire g24916;
wire II30617;
wire g10690;
wire II17705;
wire g28417;
wire g30873;
wire II18341;
wire g24855;
wire II35518;
wire g29412;
wire g11951;
wire g9626;
wire g27204;
wire g17701;
wire g5701;
wire g9019;
wire g24712;
wire g29721;
wire g23681;
wire g28218;
wire II31607;
wire II29439;
wire II32868;
wire g8169;
wire II39794;
wire g15595;
wire g4711;
wire II36153;
wire g18630;
wire g8888;
wire g25735;
wire g16127;
wire g30474;
wire II28126;
wire g16540;
wire g27993;
wire g28034;
wire g15513;
wire g28667;
wire II29386;
wire g30905;
wire g10256;
wire g16923;
wire g22708;
wire g18808;
wire g29671;
wire g19587;
wire g11725;
wire g24094;
wire g23037;
wire g26342;
wire g5635;
wire g19633;
wire g21077;
wire g17315;
wire g30978;
wire g15981;
wire g24307;
wire g11659;
wire g7545;
wire g6149;
wire g20595;
wire g23469;
wire g8311;
wire g23124;
wire g13579;
wire g28476;
wire g10228;
wire g30036;
wire g11577;
wire II29530;
wire g2636;
wire g30530;
wire g24750;
wire g24868;
wire g16943;
wire II15847;
wire g7558;
wire g26973;
wire II21208;
wire g20189;
wire g29999;
wire g8463;
wire g15998;
wire g15104;
wire g23318;
wire g5739;
wire g16029;
wire II25371;
wire g8948;
wire g11534;
wire g9811;
wire g24434;
wire g21388;
wire g27306;
wire g18964;
wire II22737;
wire gbuf168;
wire g28029;
wire g26032;
wire g7557;
wire II36476;
wire g23620;
wire II23751;
wire g27109;
wire g20949;
wire g14385;
wire g24352;
wire g30091;
wire II22745;
wire g4231;
wire g16543;
wire II39258;
wire g22940;
wire g8571;
wire g25042;
wire g19302;
wire g25299;
wire II33717;
wire g5941;
wire g26281;
wire g10315;
wire II14298;
wire g19036;
wire g11561;
wire g22758;
wire g18330;
wire g8464;
wire g11975;
wire g30379;
wire g10789;
wire g5986;
wire g5666;
wire II16289;
wire II13236;
wire II20700;
wire g30410;
wire II28913;
wire II39573;
wire II33903;
wire g22073;
wire g4696;
wire g23887;
wire g26865;
wire g24227;
wire g27284;
wire II25180;
wire g18536;
wire g29568;
wire g8530;
wire g24374;
wire g21961;
wire g28370;
wire g11860;
wire gbuf6;
wire g19505;
wire II33390;
wire g20850;
wire II28273;
wire g6054;
wire g27726;
wire II16961;
wire g22716;
wire g23462;
wire g10200;
wire g7694;
wire II20670;
wire g12134;
wire g9126;
wire g21087;
wire g24346;
wire g27137;
wire g28360;
wire g26278;
wire II16465;
wire II30281;
wire g19773;
wire g20923;
wire g11587;
wire g26915;
wire g14124;
wire II25533;
wire g28623;
wire II15590;
wire II32334;
wire g9640;
wire g28401;
wire II16827;
wire g20583;
wire g23608;
wire g27723;
wire g22639;
wire g26723;
wire g24767;
wire g21643;
wire g29819;
wire g29365;
wire g9941;
wire II36267;
wire g13649;
wire g12071;
wire g22731;
wire g4876;
wire II18223;
wire g25189;
wire g11746;
wire g29800;
wire g21080;
wire g9815;
wire g24030;
wire II21310;
wire g5089;
wire g17291;
wire g27379;
wire g24636;
wire g12207;
wire g19265;
wire g27587;
wire g17382;
wire g17233;
wire g24423;
wire gbuf16;
wire II15983;
wire II22554;
wire g18061;
wire g24801;
wire g27274;
wire g19624;
wire g20915;
wire g27552;
wire II17954;
wire g18584;
wire II40838;
wire g8473;
wire II40510;
wire g13750;
wire g27440;
wire II34665;
wire g30613;
wire g10934;
wire g4318;
wire g19084;
wire g6836;
wire II22938;
wire g24866;
wire II24689;
wire g17509;
wire g10299;
wire g12158;
wire g18105;
wire g26965;
wire g25851;
wire g15185;
wire g25982;
wire g23590;
wire g30307;
wire II36885;
wire g9159;
wire g21424;
wire g5853;
wire g29506;
wire II30776;
wire g19276;
wire II25041;
wire g30139;
wire g12066;
wire g29384;
wire g15237;
wire II23113;
wire g12762;
wire g10513;
wire g26439;
wire g30842;
wire II13974;
wire g29977;
wire g9079;
wire g27019;
wire g25206;
wire II30483;
wire g29271;
wire g27055;
wire g20916;
wire g24469;
wire g11623;
wire II14519;
wire g22020;
wire g11705;
wire g11570;
wire g9137;
wire g23067;
wire g28489;
wire g22749;
wire g27918;
wire g12333;
wire g9778;
wire II34411;
wire g14958;
wire g28914;
wire g29405;
wire g24311;
wire II20709;
wire II21830;
wire g30368;
wire g18870;
wire II17972;
wire II28476;
wire II32916;
wire II32431;
wire g11895;
wire g15207;
wire g11772;
wire II24436;
wire g27621;
wire g12829;
wire g24417;
wire g30116;
wire g25973;
wire g19349;
wire g12769;
wire g20893;
wire g18037;
wire g15572;
wire II36327;
wire g7578;
wire II30959;
wire g23092;
wire g4201;
wire g4535;
wire g16341;
wire g27767;
wire g29231;
wire g9522;
wire g24694;
wire g23493;
wire g30522;
wire g13466;
wire g26432;
wire g30867;
wire II32203;
wire g17118;
wire g29208;
wire g13439;
wire g8474;
wire g16094;
wire II25105;
wire g29533;
wire II26025;
wire g25961;
wire g26027;
wire g22059;
wire II33564;
wire g23302;
wire g16161;
wire g5688;
wire g28909;
wire g13057;
wire g24291;
wire g25484;
wire II39077;
wire II24038;
wire g29194;
wire g16135;
wire II22120;
wire II33630;
wire g10707;
wire g26591;
wire g26533;
wire g8893;
wire II20334;
wire g28085;
wire II27191;
wire g20799;
wire g3241;
wire g25764;
wire g16049;
wire g17203;
wire g28246;
wire g27223;
wire g29076;
wire g24792;
wire g15483;
wire g22609;
wire g30573;
wire g29988;
wire g25824;
wire g18883;
wire g15993;
wire g28084;
wire g18554;
wire II18485;
wire g22536;
wire g20424;
wire II20048;
wire gbuf194;
wire II16644;
wire g11548;
wire g25313;
wire II25722;
wire g27353;
wire g11969;
wire g8079;
wire II26630;
wire g28835;
wire g28931;
wire g9461;
wire g24467;
wire g29541;
wire g24268;
wire g20008;
wire g17369;
wire g6046;
wire II27705;
wire II34879;
wire g20499;
wire g21139;
wire g23764;
wire g12968;
wire g20147;
wire g20504;
wire II28318;
wire g21815;
wire g20067;
wire g8617;
wire g16286;
wire g19419;
wire g8008;
wire g5419;
wire g30787;
wire g18864;
wire g10221;
wire g13789;
wire g28708;
wire g28638;
wire g11840;
wire II15448;
wire g29728;
wire gbuf88;
wire g27087;
wire g21885;
wire g26299;
wire g26016;
wire g26643;
wire g24318;
wire g6781;
wire g19215;
wire g14657;
wire II16255;
wire g30709;
wire gbuf69;
wire g23831;
wire II41038;
wire g29374;
wire g25507;
wire g21756;
wire g7880;
wire gbuf90;
wire II25915;
wire g4891;
wire g11622;
wire II19426;
wire gbuf13;
wire II38024;
wire II30695;
wire II41126;
wire g23644;
wire II25031;
wire g11839;
wire II35461;
wire g14811;
wire g30567;
wire g23078;
wire g27080;
wire II30692;
wire g30313;
wire g28127;
wire II26898;
wire g29417;
wire g21771;
wire g10572;
wire g13060;
wire g30700;
wire II40008;
wire g25741;
wire g26052;
wire II30997;
wire g30516;
wire g23937;
wire g5905;
wire g22771;
wire g12327;
wire g29323;
wire g30910;
wire g24592;
wire g7727;
wire g16454;
wire g23722;
wire g30218;
wire g20104;
wire g22476;
wire g11481;
wire g26512;
wire II35087;
wire g22667;
wire II32146;
wire g15438;
wire g20302;
wire g18924;
wire g24161;
wire g12407;
wire g25259;
wire g26554;
wire g7152;
wire g20719;
wire g15930;
wire II21711;
wire II35741;
wire g19044;
wire g23606;
wire II28928;
wire II24493;
wire II36444;
wire II24380;
wire II26590;
wire g12058;
wire II30260;
wire g13453;
wire g21706;
wire II18623;
wire II37322;
wire g25652;
wire g24102;
wire g15753;
wire II37656;
wire II23808;
wire II38734;
wire g29524;
wire g23576;
wire g11478;
wire g11157;
wire g18933;
wire g4659;
wire g20354;
wire g10303;
wire g11468;
wire g10994;
wire II38157;
wire g8625;
wire g19714;
wire g5997;
wire g21400;
wire II19972;
wire g16481;
wire g23255;
wire g20287;
wire II39628;
wire II19787;
wire g9663;
wire g13150;
wire II15887;
wire g19257;
wire g17892;
wire g14068;
wire g12087;
wire g4652;
wire g23599;
wire g8769;
wire g16615;
wire g6026;
wire g5753;
wire g21801;
wire g14775;
wire II25138;
wire g24339;
wire g8100;
wire g26843;
wire g16591;
wire g29647;
wire II21443;
wire g30893;
wire g26624;
wire II16372;
wire g16402;
wire II18773;
wire g28673;
wire g21958;
wire g30920;
wire II19549;
wire II37638;
wire g14637;
wire g28014;
wire g9761;
wire g5235;
wire g6060;
wire II24532;
wire g20140;
wire II36702;
wire II23960;
wire II29969;
wire g19163;
wire g13580;
wire g26181;
wire g10600;
wire g18130;
wire II36307;
wire II32380;
wire g8961;
wire II28693;
wire g12118;
wire g23790;
wire g13283;
wire g5275;
wire g4495;
wire g15644;
wire II37077;
wire g27210;
wire g8546;
wire g20634;
wire II32370;
wire II25560;
wire g20432;
wire g29981;
wire g20408;
wire g6194;
wire g15452;
wire II24546;
wire II31613;
wire II21537;
wire g25025;
wire g30736;
wire g15527;
wire II23578;
wire g21650;
wire g27224;
wire g5760;
wire II31463;
wire g27563;
wire g19380;
wire g7590;
wire g8218;
wire g15612;
wire g13036;
wire II36111;
wire g8987;
wire g20714;
wire g28329;
wire g22760;
wire II22820;
wire II18356;
wire g30696;
wire g16393;
wire g6067;
wire II38434;
wire g18058;
wire II20497;
wire g15805;
wire g22297;
wire g29452;
wire II24228;
wire g10352;
wire g20401;
wire g18561;
wire II27349;
wire II26432;
wire g12507;
wire g24383;
wire g25471;
wire g29893;
wire g21379;
wire g23305;
wire II16147;
wire II26745;
wire II15372;
wire g6626;
wire II23493;
wire g12262;
wire II15271;
wire g26148;
wire g24816;
wire g22357;
wire g15717;
wire II29638;
wire g12036;
wire II37999;
wire g28852;
wire g19894;
wire g12063;
wire g24134;
wire g21278;
wire g9471;
wire g11517;
wire g29001;
wire II18518;
wire II25084;
wire g23188;
wire g30318;
wire II25459;
wire II36647;
wire g26336;
wire II40326;
wire g30548;
wire g20606;
wire II30722;
wire II15538;
wire g28767;
wire g14419;
wire II23351;
wire g13179;
wire II26624;
wire g22101;
wire g12756;
wire II25201;
wire g28645;
wire II24943;
wire g24549;
wire g22014;
wire g15491;
wire g24668;
wire g13316;
wire g22290;
wire g14176;
wire II34851;
wire g24077;
wire II21511;
wire g11684;
wire g22305;
wire g7605;
wire g29102;
wire g15407;
wire II25338;
wire g26194;
wire II24428;
wire g17191;
wire g30917;
wire g28093;
wire II18244;
wire g26482;
wire II37164;
wire g21682;
wire g17086;
wire g10387;
wire II33918;
wire g23250;
wire g16369;
wire II31622;
wire g5977;
wire g13634;
wire II19211;
wire II22946;
wire g20014;
wire g21787;
wire g5718;
wire g20443;
wire g19049;
wire II30131;
wire g27494;
wire g8360;
wire II14688;
wire g11355;
wire g5420;
wire g13527;
wire g12467;
wire g28233;
wire II32265;
wire g18446;
wire g5349;
wire II29033;
wire II21995;
wire g15080;
wire g26582;
wire g14677;
wire g11450;
wire II15873;
wire g5727;
wire g6643;
wire g11791;
wire II18238;
wire g16000;
wire g22207;
wire g4629;
wire g24215;
wire g13589;
wire g12248;
wire g27658;
wire II36650;
wire II33551;
wire g25186;
wire g23191;
wire g11580;
wire II38909;
wire II34201;
wire g17951;
wire g29787;
wire g17313;
wire g8725;
wire g30588;
wire II15893;
wire g23897;
wire II25415;
wire g25367;
wire II21755;
wire g25466;
wire g17124;
wire g24348;
wire II28087;
wire g5756;
wire g4833;
wire II37736;
wire g28791;
wire II25074;
wire g24214;
wire g15782;
wire g30199;
wire gbuf153;
wire g27111;
wire g22409;
wire g27719;
wire g9097;
wire II31742;
wire II17715;
wire g23015;
wire g25336;
wire g10150;
wire II20490;
wire g12472;
wire g24827;
wire g20255;
wire g24452;
wire g14217;
wire g5990;
wire g8841;
wire g30685;
wire g13883;
wire II38014;
wire g13602;
wire g9144;
wire g12389;
wire g27262;
wire g20295;
wire II30404;
wire g18905;
wire II18049;
wire g14719;
wire g25078;
wire g30655;
wire g22035;
wire II37587;
wire g18971;
wire g8684;
wire g10580;
wire g11990;
wire g26851;
wire g15818;
wire g17121;
wire g21003;
wire II18441;
wire g20513;
wire g20326;
wire g4398;
wire II13742;
wire g12514;
wire g7838;
wire g28263;
wire g22146;
wire g16514;
wire g11596;
wire II34719;
wire g24505;
wire g21218;
wire II36046;
wire g12296;
wire g11554;
wire g13619;
wire g12462;
wire gbuf70;
wire g27217;
wire g13342;
wire g20048;
wire g19548;
wire g4182;
wire g30003;
wire g30066;
wire g30078;
wire g30457;
wire g29379;
wire g29839;
wire g9335;
wire II21566;
wire g4000;
wire II36906;
wire g27764;
wire g27463;
wire g23439;
wire II25067;
wire g28386;
wire g28710;
wire g25245;
wire g11529;
wire II24486;
wire II27125;
wire g13122;
wire II32285;
wire g10357;
wire II28766;
wire g19819;
wire g26136;
wire g8968;
wire g10179;
wire g28666;
wire g22740;
wire II33614;
wire g30183;
wire II40739;
wire g20451;
wire g3774;
wire g15392;
wire g9907;
wire II18198;
wire II39866;
wire II20673;
wire g25170;
wire g26199;
wire II30020;
wire g15651;
wire II14525;
wire g26440;
wire II25557;
wire II38659;
wire II25624;
wire II38456;
wire II27838;
wire g4610;
wire II27352;
wire g28996;
wire II18145;
wire II36803;
wire g29214;
wire II17658;
wire g19948;
wire g10195;
wire g20999;
wire II36280;
wire g27510;
wire g17676;
wire g18062;
wire II15469;
wire II40640;
wire II40637;
wire g30692;
wire II29067;
wire g10042;
wire g24517;
wire II29629;
wire g16413;
wire g8090;
wire g27116;
wire g13431;
wire II37824;
wire g12772;
wire II25114;
wire II37095;
wire g19585;
wire II24299;
wire g7763;
wire gbuf156;
wire g10535;
wire II24156;
wire g27773;
wire g22610;
wire g16051;
wire g19781;
wire g14766;
wire II19226;
wire g15722;
wire g30357;
wire II31310;
wire g22386;
wire g5788;
wire g6293;
wire g11249;
wire g5711;
wire g29810;
wire g28871;
wire g28010;
wire II32624;
wire g5748;
wire g14244;
wire g5805;
wire II16838;
wire g5216;
wire g7352;
wire II40104;
wire g18980;
wire g24884;
wire II31526;
wire g30725;
wire g13971;
wire g14737;
wire g8537;
wire g12811;
wire II14559;
wire g10571;
wire g9785;
wire g17084;
wire II27098;
wire g20683;
wire g29477;
wire g20332;
wire g15658;
wire II22014;
wire g18973;
wire g18567;
wire g22577;
wire II23498;
wire II25710;
wire II25395;
wire II27023;
wire g16427;
wire g26706;
wire II33000;
wire g13151;
wire g6022;
wire II30847;
wire g4985;
wire g17585;
wire II14786;
wire II25781;
wire g24587;
wire g8532;
wire g8403;
wire g28261;
wire II16134;
wire g6222;
wire g13101;
wire II29881;
wire g27199;
wire g29499;
wire II20131;
wire g21005;
wire II32297;
wire g13140;
wire II34343;
wire gbuf71;
wire g4401;
wire g28256;
wire II18608;
wire g13408;
wire g9879;
wire II24326;
wire g26583;
wire g20083;
wire II29366;
wire g28077;
wire II31754;
wire II35383;
wire II25258;
wire g7604;
wire g19420;
wire g21804;
wire II15938;
wire g28882;
wire g20776;
wire II18058;
wire II33603;
wire II36780;
wire II24588;
wire g12085;
wire g7192;
wire g29844;
wire g28266;
wire II39853;
wire g29762;
wire g30941;
wire g22587;
wire II40021;
wire g22839;
wire II36087;
wire g10176;
wire g8779;
wire g17045;
wire II26571;
wire II37471;
wire g19491;
wire II23888;
wire g16679;
wire II19563;
wire g26381;
wire g13700;
wire II35809;
wire g29611;
wire g18966;
wire g12256;
wire g4421;
wire g7895;
wire g19829;
wire g19899;
wire g25375;
wire g28523;
wire g22213;
wire II21458;
wire II15505;
wire g19598;
wire g28721;
wire g29225;
wire g19498;
wire g14175;
wire gbuf217;
wire g16200;
wire g12173;
wire II32368;
wire g13846;
wire g7626;
wire g22767;
wire g16424;
wire g30369;
wire g13563;
wire II30266;
wire g30948;
wire g22132;
wire g26324;
wire g19110;
wire g13165;
wire g5694;
wire II18719;
wire g20616;
wire g18085;
wire g15556;
wire II28072;
wire g12329;
wire g19744;
wire II18142;
wire II27711;
wire g30543;
wire g23882;
wire g19836;
wire g19149;
wire II17963;
wire g30755;
wire g28671;
wire g28039;
wire g26947;
wire g20467;
wire gbuf203;
wire II18458;
wire II23065;
wire g23632;
wire g13286;
wire g17776;
wire II22064;
wire II27984;
wire g4144;
wire II35678;
wire g13819;
wire g28327;
wire II17653;
wire g23173;
wire g29430;
wire II30575;
wire II34464;
wire II22973;
wire g20878;
wire g28284;
wire g8520;
wire II37611;
wire II39264;
wire II35714;
wire g28940;
wire g13946;
wire g14883;
wire II32645;
wire g27503;
wire g28735;
wire g23673;
wire g28060;
wire II18007;
wire g15528;
wire g26853;
wire II29080;
wire g19132;
wire g9149;
wire g13736;
wire g5758;
wire g28290;
wire II33009;
wire II27264;
wire II20504;
wire II38820;
wire II21871;
wire g24390;
wire II26564;
wire II38931;
wire g23675;
wire g25389;
wire g17405;
wire g25470;
wire g24490;
wire g19554;
wire g10625;
wire II34316;
wire g20279;
wire g16240;
wire g16682;
wire g5958;
wire II34083;
wire g26747;
wire g27222;
wire g13074;
wire g9764;
wire II13194;
wire II33324;
wire g18520;
wire II31718;
wire g27259;
wire g20382;
wire g25291;
wire g29484;
wire g17304;
wire g5814;
wire g12797;
wire II16656;
wire g27515;
wire II32633;
wire g24002;
wire g22829;
wire II26679;
wire g24823;
wire g19802;
wire g15770;
wire g13953;
wire II20823;
wire II37068;
wire g25117;
wire II23377;
wire g24168;
wire II30251;
wire g17900;
wire g12883;
wire g13517;
wire g11710;
wire g28817;
wire g24997;
wire II27577;
wire g10374;
wire II26413;
wire g11886;
wire g29514;
wire g10366;
wire g9384;
wire g22586;
wire g25150;
wire g9041;
wire II15869;
wire g12979;
wire II35829;
wire g11913;
wire g6055;
wire g4266;
wire II19774;
wire II22954;
wire g26311;
wire II32946;
wire g26845;
wire g28382;
wire g23231;
wire g27400;
wire g26005;
wire g26984;
wire g11706;
wire II34159;
wire g10320;
wire II25579;
wire g19981;
wire g18974;
wire g8558;
wire g26050;
wire g9215;
wire g29284;
wire II23866;
wire g12293;
wire g29465;
wire g12786;
wire II18368;
wire g12893;
wire g29919;
wire g20507;
wire g28665;
wire g29136;
wire II31481;
wire g21334;
wire g27407;
wire II27419;
wire g26740;
wire g22091;
wire g29631;
wire g13176;
wire g7925;
wire g11870;
wire g21440;
wire gbuf60;
wire g29557;
wire g29002;
wire g16671;
wire g22157;
wire g29042;
wire g15667;
wire II24744;
wire g29322;
wire g21313;
wire g19735;
wire g28274;
wire g10471;
wire g12163;
wire II18067;
wire g13080;
wire g13108;
wire II16228;
wire g28351;
wire g21357;
wire g24580;
wire g5159;
wire II37182;
wire g27322;
wire g5396;
wire II39892;
wire g21355;
wire gbuf64;
wire g11523;
wire gbuf139;
wire g22603;
wire g7996;
wire g19290;
wire g21084;
wire g13450;
wire g8673;
wire g26447;
wire g13446;
wire g9524;
wire II32661;
wire g26593;
wire II30870;
wire g27104;
wire g27335;
wire g24969;
wire g11540;
wire g25018;
wire II22025;
wire g28460;
wire g17016;
wire g26427;
wire g25790;
wire g16626;
wire g17064;
wire II37323;
wire II28380;
wire g30241;
wire g24316;
wire II17724;
wire g7484;
wire II27992;
wire g16452;
wire g10499;
wire II14143;
wire II38348;
wire g8340;
wire g8004;
wire II18426;
wire g30305;
wire g23668;
wire g29144;
wire g12102;
wire g30676;
wire g19687;
wire II15433;
wire II22630;
wire g27031;
wire g24952;
wire II15815;
wire g24153;
wire g22921;
wire II16720;
wire g12455;
wire g28446;
wire g8489;
wire II40976;
wire II16524;
wire g19010;
wire II30188;
wire g28579;
wire II28649;
wire g26545;
wire II32491;
wire II32392;
wire g21732;
wire g30632;
wire II21595;
wire II29348;
wire g21569;
wire g10523;
wire g29792;
wire II31709;
wire g30622;
wire g9644;
wire II40173;
wire g27237;
wire g23331;
wire II29741;
wire g19734;
wire II40603;
wire g9583;
wire II39023;
wire g28150;
wire II13868;
wire g10395;
wire II29984;
wire g12023;
wire g26085;
wire g15399;
wire g10814;
wire II28248;
wire g26084;
wire g26366;
wire II38749;
wire g20809;
wire g22399;
wire g12437;
wire g29622;
wire g25821;
wire g14524;
wire II39276;
wire g24619;
wire g28032;
wire II16114;
wire II25225;
wire II32419;
wire g22675;
wire g15758;
wire g16293;
wire II28435;
wire g8525;
wire g21631;
wire g12980;
wire II36096;
wire g7830;
wire g11441;
wire II26472;
wire g12145;
wire g10726;
wire g4076;
wire II23920;
wire g21849;
wire g26417;
wire II23265;
wire g27263;
wire II39689;
wire II27134;
wire II40778;
wire II40748;
wire g21694;
wire g17093;
wire II23692;
wire g12848;
wire g6226;
wire g30329;
wire g14015;
wire g29387;
wire II25057;
wire g9808;
wire g5676;
wire g13241;
wire g25939;
wire g28289;
wire g10450;
wire g13468;
wire g20223;
wire g4225;
wire g29228;
wire II15636;
wire g23586;
wire g22241;
wire II25826;
wire g26962;
wire II24112;
wire gbuf123;
wire g15734;
wire g12515;
wire g5312;
wire g13064;
wire II24633;
wire II36728;
wire g5687;
wire g28641;
wire g11693;
wire II29004;
wire g10231;
wire g22193;
wire II21926;
wire g21045;
wire g20162;
wire g11185;
wire II22947;
wire g25190;
wire g13385;
wire II21989;
wire g10158;
wire g23246;
wire g26350;
wire g9953;
wire g25984;
wire g27443;
wire g11786;
wire g18948;
wire g24428;
wire g15243;
wire g15952;
wire g8068;
wire g19889;
wire II21337;
wire g26950;
wire g23640;
wire g10638;
wire II26651;
wire g12077;
wire g23819;
wire g26760;
wire g20120;
wire g20386;
wire II34644;
wire g29627;
wire g17560;
wire g15680;
wire g10448;
wire II39870;
wire g12548;
wire g14091;
wire g12098;
wire II35897;
wire g25969;
wire g12037;
wire g19048;
wire g9424;
wire II33885;
wire II25772;
wire g21423;
wire g19691;
wire g27003;
wire II18070;
wire g17837;
wire g19614;
wire g20910;
wire g11208;
wire II18596;
wire g18247;
wire II23679;
wire II30356;
wire II16581;
wire g20099;
wire g17281;
wire II40310;
wire g19268;
wire g5242;
wire g26844;
wire g30875;
wire g3253;
wire g26309;
wire g21544;
wire g25199;
wire g30740;
wire g23226;
wire g26451;
wire g29503;
wire II29252;
wire g13670;
wire II23371;
wire II32991;
wire g20348;
wire II21894;
wire g9790;
wire II25888;
wire g6044;
wire g17667;
wire II21979;
wire g5846;
wire II16711;
wire g24837;
wire g24242;
wire g11642;
wire g26735;
wire g29309;
wire g24905;
wire II25237;
wire g25011;
wire II21900;
wire g30059;
wire g12432;
wire g23281;
wire II30068;
wire g11810;
wire II19877;
wire II37269;
wire g26633;
wire g30747;
wire g5937;
wire g29296;
wire g4916;
wire g4954;
wire g9909;
wire g22064;
wire II23309;
wire g23240;
wire g20412;
wire g30790;
wire g20956;
wire g7635;
wire g13997;
wire II40507;
wire g29104;
wire g22979;
wire g24368;
wire g6102;
wire g17352;
wire g25543;
wire II33257;
wire g18931;
wire II39991;
wire g22696;
wire g21125;
wire II27332;
wire II23454;
wire II29841;
wire II17942;
wire II29215;
wire g28920;
wire II21629;
wire II20583;
wire g11231;
wire g22245;
wire g10518;
wire g15264;
wire g26611;
wire g26506;
wire g13237;
wire g26647;
wire g18812;
wire II21694;
wire g14797;
wire g29610;
wire g18190;
wire g20582;
wire II31940;
wire II25183;
wire g25585;
wire g21708;
wire g4451;
wire g19207;
wire g14328;
wire g5979;
wire II30218;
wire g26014;
wire g30803;
wire II36270;
wire g30377;
wire gbuf142;
wire II20828;
wire g24403;
wire II33873;
wire II18115;
wire g23555;
wire g16044;
wire g26654;
wire g30629;
wire g13092;
wire g8646;
wire II23622;
wire II27185;
wire g12558;
wire g28051;
wire g17673;
wire g7562;
wire g18024;
wire g24353;
wire g16485;
wire II39145;
wire II15771;
wire II32877;
wire II35347;
wire g24858;
wire II15466;
wire g24521;
wire g18616;
wire II34121;
wire g8703;
wire g28125;
wire g26349;
wire g16012;
wire g11643;
wire g30502;
wire g22027;
wire g20221;
wire g24249;
wire g21432;
wire g4479;
wire g18636;
wire g8651;
wire g22332;
wire II30751;
wire g13162;
wire II36987;
wire g30090;
wire II18650;
wire g16461;
wire g5914;
wire g21820;
wire g26710;
wire g16909;
wire g25932;
wire gbuf4;
wire g28295;
wire g28091;
wire II37104;
wire g19766;
wire g16100;
wire g5777;
wire g14033;
wire II13993;
wire g14221;
wire II33338;
wire g10485;
wire II14739;
wire II13947;
wire g30475;
wire II30098;
wire g28829;
wire g21025;
wire g8287;
wire II33289;
wire II15460;
wire g12486;
wire II35893;
wire II36800;
wire g9605;
wire g25958;
wire g11923;
wire g29393;
wire g30931;
wire g28161;
wire II18420;
wire g20453;
wire II25177;
wire II24144;
wire g24445;
wire g8053;
wire g16794;
wire g8497;
wire II31074;
wire g27185;
wire g22637;
wire g25224;
wire g12123;
wire g15218;
wire g10406;
wire g26302;
wire g30295;
wire g29939;
wire g20497;
wire g9869;
wire II25816;
wire g30639;
wire g11031;
wire g29363;
wire g23842;
wire g24089;
wire g21527;
wire II33558;
wire g23908;
wire g20615;
wire II23415;
wire g5936;
wire g10765;
wire g27564;
wire g27272;
wire g13256;
wire g20192;
wire g29348;
wire g21795;
wire g17269;
wire g28874;
wire II18274;
wire g23859;
wire g20754;
wire g7228;
wire II20529;
wire g30717;
wire g30317;
wire g22686;
wire g30559;
wire II26525;
wire II25120;
wire II35703;
wire g26627;
wire g12000;
wire g15866;
wire II15226;
wire II14459;
wire g11685;
wire g19745;
wire g26303;
wire g20182;
wire g12692;
wire g26773;
wire g30211;
wire g12933;
wire g23496;
wire II33542;
wire g13048;
wire g26818;
wire g19696;
wire g8555;
wire g7857;
wire g28846;
wire g25927;
wire g16477;
wire g8172;
wire II19469;
wire g8138;
wire g6512;
wire g28422;
wire g25214;
wire II27068;
wire g5379;
wire II33405;
wire II30341;
wire II16867;
wire g19313;
wire g19798;
wire g4865;
wire g23001;
wire g21060;
wire II25525;
wire g17139;
wire II21598;
wire g14529;
wire g17468;
wire g15579;
wire g19441;
wire II29154;
wire g11901;
wire g21725;
wire g21069;
wire g20757;
wire g10559;
wire g18758;
wire g30820;
wire g28319;
wire II14825;
wire g19850;
wire II38169;
wire II40907;
wire g3649;
wire g24226;
wire II16541;
wire II34105;
wire II21241;
wire g12922;
wire II30146;
wire g24131;
wire g8500;
wire g10496;
wire g15857;
wire g22902;
wire g22874;
wire II38193;
wire g27456;
wire II28962;
wire II21862;
wire g16497;
wire g21208;
wire g10114;
wire g21269;
wire g22285;
wire g4708;
wire g5186;
wire II30206;
wire g24377;
wire g20725;
wire g23267;
wire II20745;
wire g30151;
wire g27524;
wire g30710;
wire II36990;
wire g5981;
wire g22141;
wire II30642;
wire g19157;
wire g11906;
wire II16085;
wire g24058;
wire g18225;
wire g10334;
wire g20641;
wire g6310;
wire g9913;
wire II29909;
wire II20610;
wire II40272;
wire g23002;
wire g22000;
wire II18791;
wire g13182;
wire II14052;
wire g28113;
wire g29829;
wire g15912;
wire g21412;
wire II24258;
wire g23451;
wire II14596;
wire g29245;
wire g27903;
wire g16031;
wire g16987;
wire II25994;
wire g26398;
wire II32369;
wire g18258;
wire g17847;
wire g18165;
wire g7230;
wire II19539;
wire g22595;
wire g19859;
wire g21891;
wire II38175;
wire g21869;
wire g16391;
wire g24510;
wire g23773;
wire g11492;
wire g21149;
wire g13478;
wire g13238;
wire II25773;
wire II23433;
wire g9125;
wire g20308;
wire g27178;
wire g28185;
wire II19526;
wire g17408;
wire II33968;
wire II20565;
wire g30888;
wire g4821;
wire g16276;
wire g25035;
wire g11088;
wire g19024;
wire g26207;
wire II33692;
wire g13097;
wire II27071;
wire g26166;
wire g14301;
wire g7667;
wire II21452;
wire g20445;
wire II36159;
wire II15822;
wire g30601;
wire g19202;
wire II31877;
wire II14475;
wire g18555;
wire g23133;
wire g26053;
wire II36930;
wire II40958;
wire g10164;
wire g20589;
wire g16229;
wire II30317;
wire g13416;
wire g13490;
wire II37894;
wire g27318;
wire g29165;
wire g10749;
wire II39139;
wire II38810;
wire g28338;
wire g30527;
wire g7477;
wire g26409;
wire g15129;
wire g23912;
wire g27299;
wire g19389;
wire g28611;
wire g7462;
wire II39041;
wire g6048;
wire g23032;
wire g8294;
wire g23789;
wire II24132;
wire II24727;
wire g15521;
wire II36135;
wire g5035;
wire II18482;
wire II34909;
wire g15422;
wire g11021;
wire g15932;
wire g10223;
wire II38623;
wire II38187;
wire g27064;
wire g17794;
wire g19935;
wire II24764;
wire g23013;
wire II22530;
wire II29669;
wire g11551;
wire g28803;
wire g27776;
wire g7682;
wire g21245;
wire g15351;
wire g8363;
wire g21914;
wire II15499;
wire II29220;
wire g4842;
wire II35968;
wire g22277;
wire g16085;
wire g7388;
wire g23218;
wire II14715;
wire g11219;
wire g28754;
wire g25602;
wire g22592;
wire g18896;
wire g24256;
wire g30338;
wire g29940;
wire g30904;
wire g16851;
wire II39360;
wire g28209;
wire g12520;
wire II34770;
wire g8667;
wire g18916;
wire II36870;
wire g19650;
wire g26210;
wire g23628;
wire g15563;
wire g18911;
wire g30351;
wire g7842;
wire g29200;
wire g12527;
wire g11761;
wire g30569;
wire g10763;
wire II15206;
wire II28949;
wire II40487;
wire II38064;
wire II23278;
wire II37065;
wire g13551;
wire II22062;
wire g12450;
wire g26875;
wire g18155;
wire g30771;
wire g24080;
wire g17180;
wire g13353;
wire g29159;
wire II24382;
wire g18955;
wire II37808;
wire g25136;
wire g18537;
wire g10082;
wire g10105;
wire g19591;
wire g21740;
wire g15305;
wire g23564;
wire g26521;
wire g27817;
wire II37771;
wire g6130;
wire II32985;
wire g20967;
wire g9326;
wire g20989;
wire II29915;
wire g28176;
wire II39367;
wire g23270;
wire II18758;
wire g11240;
wire g29319;
wire II35360;
wire II16605;
wire g29023;
wire g23825;
wire g4769;
wire II36633;
wire g13197;
wire g15495;
wire g16266;
wire g23353;
wire II14568;
wire g13611;
wire g23763;
wire g30383;
wire g20419;
wire II26561;
wire g23257;
wire II31664;
wire g8132;
wire g16924;
wire g20708;
wire II23530;
wire g17791;
wire g4093;
wire II41093;
wire g9119;
wire g13497;
wire II17783;
wire II21045;
wire g29189;
wire g24148;
wire g24474;
wire II21551;
wire g25168;
wire g23275;
wire g28790;
wire II14628;
wire II15626;
wire g23481;
wire g13906;
wire g28146;
wire g18839;
wire g11079;
wire g23862;
wire g18938;
wire g4800;
wire g8622;
wire g10055;
wire g26573;
wire g29099;
wire g22106;
wire g17570;
wire g21154;
wire g28221;
wire g24289;
wire g30287;
wire g11856;
wire g10587;
wire g28402;
wire g7342;
wire g4436;
wire g4509;
wire g29350;
wire g11847;
wire g27709;
wire II40808;
wire g5623;
wire II15169;
wire g22402;
wire II22593;
wire g19630;
wire II25618;
wire II25358;
wire II39809;
wire g9928;
wire g24556;
wire g21098;
wire II18635;
wire g11536;
wire g10049;
wire g16310;
wire g23458;
wire II24400;
wire g12067;
wire g15470;
wire g24385;
wire g8256;
wire g23692;
wire g27786;
wire g10723;
wire g30645;
wire g12860;
wire g12366;
wire II39392;
wire II31856;
wire g25818;
wire II31213;
wire g14753;
wire II29036;
wire II18028;
wire g25269;
wire g26717;
wire II23227;
wire g21300;
wire g23784;
wire II37644;
wire II13089;
wire g27949;
wire II18235;
wire g27025;
wire g19379;
wire g24238;
wire II34385;
wire g10652;
wire II37426;
wire g27038;
wire II32520;
wire II18659;
wire g30788;
wire g20228;
wire g28088;
wire g30220;
wire g16185;
wire g19220;
wire g30707;
wire g25834;
wire II24133;
wire g26615;
wire g17877;
wire g16109;
wire g26901;
wire II22475;
wire g15092;
wire g5406;
wire II22893;
wire g28760;
wire II32679;
wire II27235;
wire II34758;
wire g7483;
wire g10847;
wire g8566;
wire g10842;
wire g22726;
wire II29378;
wire g25357;
wire g23509;
wire g24230;
wire g19729;
wire g12006;
wire g25159;
wire gbuf212;
wire II41111;
wire II27761;
wire g29090;
wire II30501;
wire II22694;
wire II24982;
wire g20318;
wire g22293;
wire g8921;
wire II36530;
wire g30167;
wire g14414;
wire g19210;
wire g30585;
wire g27674;
wire g30375;
wire II25204;
wire g11612;
wire II29930;
wire II18647;
wire g6568;
wire g21880;
wire II21377;
wire g6063;
wire g23117;
wire g25087;
wire II25567;
wire g15858;
wire II31508;
wire g30925;
wire II30669;
wire g29215;
wire g12060;
wire g17194;
wire II23323;
wire g5992;
wire II22566;
wire g20550;
wire II18614;
wire g17567;
wire II18064;
wire g19330;
wire II16915;
wire II23581;
wire g13246;
wire g8850;
wire g29126;
wire g12510;
wire g26456;
wire g21299;
wire gbuf44;
wire II25751;
wire g20559;
wire II21508;
wire g20603;
wire g18486;
wire gbuf186;
wire g6431;
wire II35915;
wire g25744;
wire g28655;
wire g11512;
wire II30368;
wire II27958;
wire g10340;
wire II30071;
wire II28084;
wire g27846;
wire g10456;
wire II37086;
wire II26910;
wire II25683;
wire g24113;
wire g20476;
wire g19197;
wire g9438;
wire g15824;
wire g24279;
wire g29789;
wire II23524;
wire g26317;
wire g23794;
wire II36615;
wire g21888;
wire g29984;
wire g10353;
wire g26190;
wire II27868;
wire II23879;
wire II17627;
wire g30580;
wire g25476;
wire g13078;
wire g29543;
wire g5823;
wire g19138;
wire g12973;
wire g25334;
wire g20568;
wire gbuf36;
wire g16473;
wire g26754;
wire g29490;
wire g16860;
wire g22835;
wire II24093;
wire II29572;
wire g8357;
wire g25384;
wire g29459;
wire g12999;
wire g25254;
wire II23329;
wire g5230;
wire II28609;
wire g22303;
wire g4772;
wire g22078;
wire II25047;
wire g19117;
wire II37194;
wire g17207;
wire g15507;
wire gbuf111;
wire II28219;
wire g11494;
wire II24619;
wire g27578;
wire g26623;
wire g9755;
wire g20144;
wire g14580;
wire g22233;
wire g16090;
wire g19169;
wire II36957;
wire g18828;
wire g30962;
wire g25957;
wire g29757;
wire g17617;
wire g20519;
wire g16071;
wire II24148;
wire II13604;
wire g5955;
wire II34002;
wire g7146;
wire g5850;
wire g26049;
wire II31005;
wire II29622;
wire g25331;
wire g12272;
wire g4366;
wire g18174;
wire g18189;
wire g19620;
wire g27201;
wire g18669;
wire g7989;
wire g16112;
wire g20866;
wire II29966;
wire g22882;
wire II31898;
wire g19663;
wire g30005;
wire g21033;
wire g30027;
wire g8541;
wire II29104;
wire g20329;
wire g12644;
wire g15321;
wire II22869;
wire g21655;
wire g9527;
wire g23832;
wire g4818;
wire g8689;
wire II17100;
wire g21487;
wire g10304;
wire gbuf56;
wire II40628;
wire II22284;
wire II36221;
wire g24414;
wire g30659;
wire II16034;
wire g11583;
wire gbuf9;
wire g17200;
wire g30501;
wire g27714;
wire g13524;
wire II26892;
wire g18231;
wire II34254;
wire g30652;
wire g24282;
wire g12266;
wire II23794;
wire g16069;
wire II25898;
wire II22741;
wire g8621;
wire II25913;
wire II23959;
wire g21686;
wire II17701;
wire g19484;
wire g5546;
wire g25462;
wire g13535;
wire II18497;
wire g20975;
wire g23198;
wire g27763;
wire g27495;
wire g27465;
wire g18922;
wire g19170;
wire g5767;
wire g29912;
wire g19064;
wire II24063;
wire g9074;
wire g9889;
wire g21187;
wire g6281;
wire g30409;
wire g10888;
wire g16401;
wire II22855;
wire II38905;
wire g24509;
wire g5418;
wire g27213;
wire g17099;
wire g24502;
wire g20896;
wire g17115;
wire g11843;
wire g15840;
wire g21845;
wire g22003;
wire g11593;
wire g25364;
wire II32955;
wire g13817;
wire g17862;
wire II22690;
wire g20304;
wire g12130;
wire g5343;
wire g30464;
wire II23436;
wire g27630;
wire g13155;
wire g20899;
wire g5338;
wire g15817;
wire g11525;
wire g28932;
wire g28692;
wire g28394;
wire g23253;
wire g27076;
wire g4314;
wire II25463;
wire g5750;
wire g20321;
wire g9933;
wire g14213;
wire g9263;
wire g26384;
wire g22738;
wire g20291;
wire II36382;
wire g19700;
wire g24682;
wire g18091;
wire g19927;
wire g13573;
wire g27394;
wire II16566;
wire g25527;
wire g29564;
wire g26310;
wire g10172;
wire II16261;
wire g19763;
wire g6021;
wire g30009;
wire II39032;
wire g16288;
wire II30086;
wire II15523;
wire g12901;
wire g26437;
wire g27627;
wire II21271;
wire g27560;
wire g11944;
wire II30176;
wire g15389;
wire g24217;
wire gbuf77;
wire g12991;
wire g28501;
wire g30681;
wire g30784;
wire g22649;
wire II24338;
wire g11729;
wire g25174;
wire g27381;
wire g25328;
wire g18407;
wire g26881;
wire g27656;
wire g3969;
wire g29054;
wire g19382;
wire II24307;
wire II19844;
wire g13854;
wire g13886;
wire g21477;
wire II19401;
wire II36644;
wire g23767;
wire g10805;
wire II39127;
wire II30005;
wire g10144;
wire g9287;
wire g12336;
wire g11775;
wire g8821;
wire II38854;
wire g11964;
wire g23428;
wire g29400;
wire g8826;
wire g5070;
wire g5857;
wire II22551;
wire g13494;
wire II37026;
wire g4851;
wire g17237;
wire g27720;
wire g10869;
wire g22644;
wire g24397;
wire g27010;
wire II25442;
wire g29684;
wire g26075;
wire g26251;
wire II33900;
wire II24062;
wire II18205;
wire g27357;
wire g7670;
wire g22619;
wire g27250;
wire II24684;
wire g13296;
wire g7426;
wire II30790;
wire g26822;
wire g15592;
wire g5741;
wire g29580;
wire g21262;
wire g22852;
wire g28706;
wire II21661;
wire g20579;
wire g21371;
wire g13266;
wire g19475;
wire II29900;
wire g23874;
wire g15838;
wire g8670;
wire g8718;
wire g15624;
wire g29700;
wire II31838;
wire II36903;
wire II35940;
wire g28906;
wire g12392;
wire gbuf216;
wire g13838;
wire g20428;
wire II14775;
wire II17819;
wire g18492;
wire II32248;
wire g9310;
wire g17493;
wire g19017;
wire g11720;
wire g9895;
wire g22473;
wire g10414;
wire II23171;
wire II36999;
wire g17397;
wire II13122;
wire II39873;
wire II38466;
wire g15585;
wire g29299;
wire gbuf199;
wire g27584;
wire g4335;
wire g5061;
wire g5923;
wire g9091;
wire II21560;
wire g11961;
wire g24121;
wire g9487;
wire g12443;
wire g19029;
wire g27684;
wire II19582;
wire g28173;
wire g9795;
wire g15030;
wire g27581;
wire g23745;
wire II36539;
wire II20832;
wire g25185;
wire g7566;
wire II17957;
wire g24543;
wire g13131;
wire II21825;
wire g8562;
wire g23666;
wire g29265;
wire g19904;
wire II26461;
wire g27914;
wire g16137;
wire g26023;
wire II33683;
wire g16594;
wire g8449;
wire g17591;
wire II24751;
wire g20840;
wire g23263;
wire II13092;
wire II28247;
wire g17111;
wire II38539;
wire II27621;
wire g13275;
wire II25015;
wire II16744;
wire g25283;
wire II14951;
wire g11671;
wire II31700;
wire II33168;
wire II24602;
wire g19887;
wire g18935;
wire II40588;
wire g29725;
wire g18128;
wire g25310;
wire g28741;
wire II17673;
wire g10263;
wire g5703;
wire g16056;
wire g15737;
wire g29656;
wire g24863;
wire g20993;
wire II22726;
wire II19360;
wire II16556;
wire g18419;
wire g4006;
wire II16486;
wire g12109;
wire g5642;
wire g17216;
wire g26371;
wire g13608;
wire g11835;
wire g19183;
wire II18801;
wire g30688;
wire g9098;
wire II21569;
wire g11628;
wire II36447;
wire g18060;
wire g17503;
wire II16870;
wire g10252;
wire g27164;
wire II21855;
wire II14848;
wire II34812;
wire g28169;
wire g4430;
wire g8783;
wire g22747;
wire g27085;
wire g18474;
wire g24539;
wire g8711;
wire g27276;
wire g21811;
wire II16059;
wire II41035;
wire g22706;
wire g22663;
wire II26028;
wire g19307;
wire g26174;
wire g19184;
wire g28702;
wire g10988;
wire g26588;
wire g24084;
wire II29055;
wire g8762;
wire II15191;
wire g9183;
wire g7224;
wire II39348;
wire g23357;
wire g11407;
wire g23799;
wire II25904;
wire g28486;
wire g9870;
wire g12765;
wire II20324;
wire g18007;
wire g10297;
wire g17189;
wire II31043;
wire II21658;
wire g24105;
wire g28745;
wire g15853;
wire g29530;
wire g24035;
wire g4609;
wire II16958;
wire g23041;
wire g5976;
wire g17162;
wire g21906;
wire g19667;
wire II35458;
wire g17948;
wire g21824;
wire gbuf18;
wire g20938;
wire g20947;
wire g10307;
wire g20177;
wire g29690;
wire g19350;
wire g24260;
wire g21374;
wire g8602;
wire g24295;
wire II27365;
wire g12053;
wire g24547;
wire g4205;
wire II22988;
wire g20563;
wire g27972;
wire g24399;
wire g21950;
wire g25243;
wire g5201;
wire g12436;
wire II19823;
wire g19675;
wire g4558;
wire II25171;
wire II25790;
wire g18121;
wire II39647;
wire g26969;
wire g22009;
wire g13620;
wire g20593;
wire g27091;
wire g27831;
wire g13457;
wire II21923;
wire II20022;
wire II40233;
wire g9120;
wire g24597;
wire g30851;
wire g19679;
wire g24333;
wire g24220;
wire g23325;
wire II40676;
wire g26595;
wire g25951;
wire g24054;
wire g25142;
wire II40459;
wire g25182;
wire g30865;
wire g29450;
wire g17992;
wire II32659;
wire g19815;
wire II33427;
wire g20351;
wire g14746;
wire g22548;
wire g11852;
wire g4783;
wire g23020;
wire g23208;
wire g19532;
wire II32452;
wire II32615;
wire g16132;
wire g11996;
wire II31775;
wire g12106;
wire g17425;
wire g25979;
wire g22032;
wire g3239;
wire g17454;
wire II18626;
wire II33894;
wire g19246;
wire g30938;
wire II34306;
wire g21338;
wire g23372;
wire g17062;
wire II30994;
wire g18276;
wire II29023;
wire II38405;
wire g16221;
wire II37313;
wire g4575;
wire g28159;
wire II36776;
wire II40221;
wire g25431;
wire g9649;
wire g20135;
wire g18328;
wire g21121;
wire g4512;
wire II28956;
wire g29380;
wire g19059;
wire II33411;
wire g22557;
wire II29426;
wire g24871;
wire g5908;
wire gbuf110;
wire g28049;
wire g8510;
wire g25784;
wire g29065;
wire g4922;
wire g27760;
wire g12187;
wire g11730;
wire g29653;
wire g27662;
wire g27157;
wire II39418;
wire g24945;
wire g7520;
wire g26802;
wire g27043;
wire II25510;
wire II34140;
wire g19095;
wire g10464;
wire g19431;
wire g18569;
wire g28774;
wire II41064;
wire g24439;
wire g16197;
wire g8901;
wire g10895;
wire II15843;
wire g11708;
wire g21947;
wire g11955;
wire g24974;
wire g26009;
wire II34535;
wire g4882;
wire II18557;
wire g22900;
wire g20284;
wire g23312;
wire II36772;
wire g21404;
wire g22152;
wire g19237;
wire II25132;
wire II34473;
wire g17500;
wire g17485;
wire g11972;
wire g30227;
wire g12539;
wire g30301;
wire II20444;
wire II24353;
wire g19603;
wire g7263;
wire II16590;
wire g29562;
wire II19624;
wire g30494;
wire II31082;
wire II24702;
wire II34044;
wire g15257;
wire g12044;
wire g10124;
wire g26038;
wire g8965;
wire II26154;
wire g20052;
wire g25860;
wire g20536;
wire g17914;
wire g23467;
wire g12379;
wire g16602;
wire II21012;
wire g6901;
wire II19587;
wire II16517;
wire g27309;
wire II23317;
wire g18787;
wire g5794;
wire g24387;
wire g9290;
wire II40820;
wire g29176;
wire g29642;
wire g24306;
wire g23601;
wire g8699;
wire g29354;
wire II14802;
wire g13227;
wire g28122;
wire g23626;
wire g26231;
wire II35946;
wire g28026;
wire g17782;
wire g8486;
wire g9022;
wire g26332;
wire g17510;
wire g11500;
wire g19936;
wire g30829;
wire g8861;
wire II15830;
wire g24762;
wire g15870;
wire g27208;
wire g24073;
wire g19502;
wire g15599;
wire II15313;
wire g28090;
wire g15710;
wire g21105;
wire g23955;
wire g4714;
wire II31568;
wire g21439;
wire g27858;
wire g24937;
wire g4677;
wire g9273;
wire g30547;
wire II16681;
wire g29964;
wire g12698;
wire II16598;
wire g23294;
wire II20100;
wire II19377;
wire g18583;
wire g30348;
wire g12180;
wire g11531;
wire II32604;
wire II32973;
wire g27538;
wire II20805;
wire g4752;
wire g27247;
wire g20218;
wire g30765;
wire g29184;
wire g11572;
wire II34677;
wire g20952;
wire II15580;
wire II15975;
wire g27728;
wire g24379;
wire g26934;
wire II32356;
wire II28068;
wire II36473;
wire g29539;
wire g13051;
wire g28435;
wire II38053;
wire g27326;
wire g27489;
wire g8107;
wire g9777;
wire g13304;
wire g5988;
wire g23870;
wire gbuf53;
wire g28270;
wire g16217;
wire II34964;
wire g20270;
wire g12113;
wire g21116;
wire g23400;
wire g5667;
wire II39767;
wire g28528;
wire g24566;
wire g21955;
wire g24320;
wire g12816;
wire g23571;
wire g18390;
wire g29152;
wire g17607;
wire g25161;
wire g27963;
wire g9000;
wire II40718;
wire g7613;
wire g19323;
wire II24544;
wire g27304;
wire g26977;
wire II21351;
wire II34168;
wire g5018;
wire II40291;
wire g18101;
wire g27267;
wire II15961;
wire g21017;
wire g28473;
wire g23048;
wire g21858;
wire g25040;
wire II37596;
wire g4684;
wire g21136;
wire g25201;
wire g9904;
wire II34740;
wire g16845;
wire II16021;
wire II23570;
wire g4386;
wire g5292;
wire g6115;
wire g7577;
wire g23407;
wire II25506;
wire g20572;
wire II31266;
wire g17321;
wire g26650;
wire II25881;
wire g28660;
wire II33617;
wire g12875;
wire g21973;
wire g28407;
wire g18690;
wire g11017;
wire g18908;
wire II29307;
wire g11930;
wire II25761;
wire II17922;
wire II18124;
wire II32687;
wire g26861;
wire II39577;
wire g17691;
wire g13030;
wire g27077;
wire g4736;
wire g20090;
wire g18804;
wire g16009;
wire g27280;
wire II32310;
wire g9634;
wire g16469;
wire II28181;
wire g20064;
wire g30832;
wire II23895;
wire II37410;
wire II17904;
wire g30393;
wire g21666;
wire II19608;
wire g21073;
wire g27931;
wire g19810;
wire g29735;
wire g8460;
wire g10259;
wire II20646;
wire g30973;
wire II37071;
wire g25021;
wire g20344;
wire g13786;
wire II33915;
wire II39939;
wire g19570;
wire II29320;
wire g12214;
wire g6033;
wire g17632;
wire g29828;
wire II13179;
wire g5872;
wire II19452;
wire g25309;
wire g29865;
wire g24965;
wire g24783;
wire g28910;
wire II30212;
wire g5969;
wire II35872;
wire gbuf143;
wire II24512;
wire g30033;
wire g26666;
wire g20984;
wire g27072;
wire g5773;
wire II39384;
wire g13645;
wire g4110;
wire g11898;
wire g8129;
wire g26501;
wire g30794;
wire g15204;
wire II32539;
wire g21326;
wire g26709;
wire g15769;
wire g8509;
wire g29927;
wire g20461;
wire g10927;
wire II38940;
wire g28193;
wire g15173;
wire II23676;
wire g13128;
wire g22184;
wire II38947;
wire g13009;
wire g22312;
wire g29193;
wire g16655;
wire II39249;
wire g26048;
wire g30485;
wire g20490;
wire g17707;
wire g23056;
wire g28714;
wire II28728;
wire g7553;
wire g24496;
wire II16182;
wire g16027;
wire g22089;
wire g7554;
wire g25049;
wire g9134;
wire II31544;
wire g7834;
wire II24251;
wire g22039;
wire II36454;
wire g25195;
wire g26727;
wire II24265;
wire g13293;
wire g21419;
wire g10991;
wire g11819;
wire g25493;
wire g11828;
wire II17916;
wire g30817;
wire g25562;
wire g19910;
wire g17577;
wire g28042;
wire g20111;
wire II16231;
wire II23689;
wire II20479;
wire II29229;
wire g13002;
wire g13112;
wire II35542;
wire g22493;
wire g10155;
wire II26532;
wire g29705;
wire g15675;
wire g16739;
wire g11808;
wire II23682;
wire II16215;
wire g26276;
wire g18429;
wire II24055;
wire g13272;
wire II13987;
wire g26263;
wire II15392;
wire II31949;
wire g21982;
wire II17898;
wire g5638;
wire II25700;
wire II15490;
wire II39886;
wire g28213;
wire g25356;
wire g22500;
wire g20440;
wire g27711;
wire g16997;
wire g22658;
wire g20655;
wire g10662;
wire g25267;
wire g20391;
wire g18851;
wire g16346;
wire g10849;
wire g21533;
wire g21197;
wire g27793;
wire g18901;
wire g30254;
wire g21091;
wire g21498;
wire II29475;
wire g21989;
wire g15022;
wire g24873;
wire II29942;
wire II25741;
wire g5881;
wire g7963;
wire g14332;
wire g30732;
wire g22308;
wire g12546;
wire g8304;
wire g19333;
wire g25518;
wire II34990;
wire g25068;
wire II30398;
wire g13541;
wire g8658;
wire g18858;
wire II14134;
wire g22118;
wire II19813;
wire g30898;
wire g3249;
wire II18587;
wire II14704;
wire g10506;
wire g25911;
wire II40937;
wire g16586;
wire g19189;
wire g8431;
wire II31274;
wire g25054;
wire g16607;
wire g26354;
wire II40862;
wire II16854;
wire g23712;
wire g22797;
wire g23639;
wire g30870;
wire II24641;
wire g29777;
wire g3994;
wire II31829;
wire II34162;
wire II31505;
wire g29772;
wire II18780;
wire g30739;
wire g18969;
wire II41129;
wire g30250;
wire g21055;
wire g24849;
wire g15404;
wire g5889;
wire II28206;
wire g12711;
wire g23128;
wire g23116;
wire g12013;
wire g22044;
wire II30493;
wire II31673;
wire II37842;
wire g20123;
wire g27926;
wire g30128;
wire g14551;
wire g6898;
wire g10224;
wire g6441;
wire II33485;
wire g11744;
wire g13250;
wire II39240;
wire g5945;
wire g18764;
wire g26073;
wire g12776;
wire g13345;
wire II37238;
wire g23855;
wire g12288;
wire g20211;
wire g28717;
wire II22044;
wire g4973;
wire II36042;
wire II34836;
wire g28497;
wire g24366;
wire g11499;
wire g29995;
wire g13205;
wire g19777;
wire g5431;
wire g29445;
wire g22270;
wire g20763;
wire g4405;
wire II19119;
wire II31595;
wire II20310;
wire II24520;
wire g23293;
wire g29013;
wire g26565;
wire g19873;
wire II25768;
wire g28688;
wire g12916;
wire gbuf109;
wire g29713;
wire II29451;
wire g4779;
wire g16337;
wire g16554;
wire g28238;
wire II37502;
wire g12234;
wire II36560;
wire g7518;
wire g19862;
wire g30886;
wire g29149;
wire g19219;
wire g4020;
wire g25885;
wire g17537;
wire g22237;
wire g11544;
wire II36510;
wire g10598;
wire g28813;
wire g30553;
wire g21381;
wire g23744;
wire g28002;
wire g21342;
wire II40604;
wire g23737;
wire g30896;
wire g30278;
wire II33440;
wire g19141;
wire g19639;
wire g7142;
wire g7973;
wire g22672;
wire g14352;
wire g30914;
wire g19504;
wire g10385;
wire g4731;
wire II23192;
wire g29806;
wire g30404;
wire g12530;
wire g6083;
wire g20626;
wire II15896;
wire II21534;
wire g27404;
wire II36945;
wire g19717;
wire g25454;
wire II21354;
wire g22679;
wire g10961;
wire II35780;
wire g18466;
wire II16763;
wire g28089;
wire g7488;
wire II36542;
wire g30449;
wire g25496;
wire g16971;
wire g29944;
wire g25628;
wire g5030;
wire II17825;
wire g11170;
wire g28796;
wire g12965;
wire II34749;
wire g14976;
wire g14478;
wire g8897;
wire g12343;
wire g28231;
wire II33463;
wire g17653;
wire g10008;
wire II27375;
wire II16098;
wire g15996;
wire gbuf102;
wire II29600;
wire g11696;
wire g30435;
wire g14904;
wire II40453;
wire g13023;
wire g18374;
wire g23618;
wire g22203;
wire g25028;
wire g8836;
wire g10604;
wire g16180;
wire g4194;
wire g5865;
wire II18034;
wire g13485;
wire g18013;
wire g17000;
wire g27346;
wire g27603;
wire g11020;
wire II32500;
wire g30903;
wire g29427;
wire g24277;
wire II27035;
wire g26784;
wire g10526;
wire g6980;
wire g27123;
wire g25260;
wire g29440;
wire g13504;
wire gbuf138;
wire g16126;
wire g18353;
wire II35467;
wire g13321;
wire II38510;
wire g26698;
wire II38223;
wire g18450;
wire g14402;
wire II14017;
wire II26494;
wire II19905;
wire g17968;
wire II35711;
wire g17333;
wire g28698;
wire g22842;
wire g28304;
wire g22626;
wire g27190;
wire II20852;
wire g22801;
wire g16383;
wire g7345;
wire II25150;
wire g6082;
wire g30959;
wire II23257;
wire II32556;
wire g26056;
wire g30122;
wire g6672;
wire II18247;
wire g29256;
wire II19611;
wire II28978;
wire g29198;
wire g23914;
wire g8394;
wire g26110;
wire g7915;
wire g12742;
wire g19033;
wire g22444;
wire g30985;
wire g21857;
wire II36789;
wire II29046;
wire g8224;
wire II24717;
wire II31141;
wire g29333;
wire g24177;
wire II40793;
wire g11135;
wire g21622;
wire II25660;
wire g25487;
wire g11095;
wire g4338;
wire g30666;
wire g12532;
wire II13433;
wire g20480;
wire g10370;
wire g11917;
wire g28341;
wire II31934;
wire g24717;
wire g13119;
wire II29897;
wire g25063;
wire g19177;
wire g5831;
wire g14007;
wire g23717;
wire g9277;
wire II35064;
wire g11508;
wire g21217;
wire g19301;
wire II26429;
wire II35500;
wire g30578;
wire g15441;
wire g18795;
wire g19549;
wire g28635;
wire g18855;
wire g16578;
wire g30261;
wire g8253;
wire g26557;
wire g22145;
wire II28272;
wire II41024;
wire g27060;
wire g26011;
wire II31766;
wire g29481;
wire II23830;
wire g12315;
wire g20503;
wire g22028;
wire gbuf68;
wire g23533;
wire g13454;
wire II36271;
wire g9286;
wire g28245;
wire g10868;
wire g30667;
wire II27739;
wire g25256;
wire II30095;
wire g9078;
wire g21350;
wire g24324;
wire II32432;
wire g4743;
wire II23839;
wire g20363;
wire g8452;
wire g19346;
wire g24571;
wire g23023;
wire II17297;
wire g22709;
wire II29052;
wire II40940;
wire II30326;
wire g18754;
wire g9520;
wire g10013;
wire g14626;
wire g30523;
wire II20664;
wire g25014;
wire g14438;
wire g15360;
wire g10324;
wire II16306;
wire g25582;
wire II39835;
wire g16160;
wire g30088;
wire II26182;
wire II40573;
wire g12354;
wire II39234;
wire g29439;
wire gbuf135;
wire II34091;
wire II29265;
wire g18200;
wire g18895;
wire g12892;
wire g25825;
wire g30872;
wire II17599;
wire g30340;
wire II31181;
wire g23107;
wire g12082;
wire g28278;
wire g20095;
wire g30967;
wire g8872;
wire II16735;
wire g15754;
wire g26464;
wire g23727;
wire g13081;
wire II14612;
wire II23729;
wire g19355;
wire g25248;
wire g29816;
wire g17645;
wire g12033;
wire g12279;
wire g17989;
wire g5173;
wire g29922;
wire g25606;
wire g29987;
wire g20421;
wire II25144;
wire II17692;
wire g10391;
wire g9227;
wire g28937;
wire g27275;
wire g26422;
wire g13442;
wire II40688;
wire II21262;
wire g11132;
wire g18689;
wire g30053;
wire II22578;
wire g13319;
wire g8869;
wire II27549;
wire g24292;
wire II39142;
wire g26223;
wire g21341;
wire g17496;
wire g4202;
wire II38863;
wire II33003;
wire g24771;
wire g10064;
wire g29229;
wire g9892;
wire g26744;
wire g23669;
wire II31472;
wire II24030;
wire g16520;
wire g22986;
wire g22920;
wire g15806;
wire II20628;
wire g25767;
wire g15151;
wire II35906;
wire g19953;
wire g6221;
wire g27311;
wire g27168;
wire g19739;
wire g12247;
wire g28333;
wire g21161;
wire g8724;
wire g30564;
wire g25352;
wire g15606;
wire g12094;
wire g8344;
wire II38217;
wire g5122;
wire g25899;
wire II16273;
wire II33424;
wire g11056;
wire g12149;
wire g30726;
wire g10423;
wire II22953;
wire g13265;
wire g29976;
wire II34051;
wire II29987;
wire II35533;
wire g16572;
wire g27678;
wire g29623;
wire g23542;
wire g6068;
wire g19563;
wire g26680;
wire II40892;
wire g20972;
wire g8156;
wire g5678;
wire II19429;
wire g17973;
wire g17594;
wire II31487;
wire g30900;
wire g18383;
wire g18207;
wire II24273;
wire g19618;
wire g10584;
wire g21184;
wire g13872;
wire II36075;
wire II38235;
wire II40727;
wire g12984;
wire II40859;
wire g26764;
wire g13056;
wire g3242;
wire g28463;
wire II36551;
wire II32608;
wire g23472;
wire II36347;
wire g25058;
wire II14030;
wire g27478;
wire II20451;
wire II24373;
wire II24453;
wire g5801;
wire g6574;
wire g28851;
wire g9523;
wire g8952;
wire II14306;
wire g18932;
wire g22102;
wire g6040;
wire II36724;
wire g23549;
wire g11782;
wire g21174;
wire g15949;
wire g4517;
wire g19738;
wire g28616;
wire g20914;
wire II24290;
wire II40745;
wire g21722;
wire g28646;
wire g13764;
wire g19411;
wire g18106;
wire g4322;
wire II28497;
wire II25819;
wire g19913;
wire II30197;
wire g23898;
wire g27998;
wire g26966;
wire g9106;
wire II33265;
wire II33316;
wire g12027;
wire II35369;
wire g22805;
wire g29383;
wire II29556;
wire g23494;
wire g27008;
wire g27396;
wire g23775;
wire g23256;
wire g21818;
wire II23028;
wire II28003;
wire g13549;
wire g23227;
wire g7742;
wire g8793;
wire g17166;
wire g30451;
wire g8574;
wire g11787;
wire g25936;
wire g25353;
wire g20986;
wire g18053;
wire II30716;
wire g24637;
wire II16238;
wire g15095;
wire g10298;
wire g29796;
wire g22127;
wire g8438;
wire g23220;
wire II29090;
wire g17243;
wire g23968;
wire g21540;
wire II23769;
wire II34647;
wire g23320;
wire II23114;
wire g28468;
wire gbuf127;
wire II30263;
wire II18289;
wire g21635;
wire g11569;
wire g23154;
wire g11562;
wire II37712;
wire g12844;
wire II13977;
wire II30713;
wire g20124;
wire II20844;
wire g19264;
wire g22401;
wire g19713;
wire g12201;
wire II26947;
wire g30673;
wire g24424;
wire g23641;
wire g29676;
wire g5428;
wire g14829;
wire II34725;
wire II15620;
wire g11836;
wire II36032;
wire g19895;
wire g11848;
wire g5715;
wire g14559;
wire g24210;
wire g7083;
wire g14837;
wire g7899;
wire g12388;
wire g19294;
wire g27112;
wire II32345;
wire g18431;
wire II34854;
wire g17633;
wire g24038;
wire g5654;
wire II37626;
wire II13224;
wire g7336;
wire II26311;
wire g28126;
wire g7348;
wire g17457;
wire g15293;
wire II31011;
wire g19805;
wire g21964;
wire g22614;
wire g26195;
wire II20676;
wire II26993;
wire g12974;
wire g19162;
wire g9044;
wire g28438;
wire gbuf152;
wire g11528;
wire II30125;
wire g20512;
wire II26334;
wire g25171;
wire g12473;
wire g13790;
wire g8775;
wire g13037;
wire g21774;
wire g11760;
wire g21873;
wire II32284;
wire g13633;
wire II23326;
wire g22622;
wire II37158;
wire II17828;
wire g30776;
wire g16421;
wire II25588;
wire g21036;
wire g23166;
wire g11606;
wire g30462;
wire g12176;
wire g24244;
wire g21677;
wire g26126;
wire gbuf146;
wire II27173;
wire g14214;
wire II36213;
wire g25394;
wire II26354;
wire g17300;
wire g11189;
wire g18319;
wire II35957;
wire g12089;
wire II31000;
wire g16529;
wire g28225;
wire II36951;
wire g7901;
wire g4346;
wire II19771;
wire g12482;
wire g16048;
wire g19092;
wire II23125;
wire II20320;
wire g16416;
wire II23142;
wire g8407;
wire II39261;
wire g11663;
wire II31823;
wire g28728;
wire II16832;
wire g26243;
wire g30934;
wire g13598;
wire g26831;
wire II39044;
wire II31805;
wire II23981;
wire II28341;
wire g22232;
wire II19573;
wire II36924;
wire g24481;
wire II40468;
wire II38502;
wire g20448;
wire g15844;
wire g8366;
wire g9058;
wire II39136;
wire g8056;
wire g17081;
wire g27798;
wire g17310;
wire II30008;
wire g29401;
wire g16142;
wire g22573;
wire g24528;
wire g24755;
wire II23386;
wire II40769;
wire g25178;
wire g17514;
wire g29472;
wire g11986;
wire g27227;
wire II29996;
wire g23157;
wire g17624;
wire II15472;
wire g26159;
wire g23095;
wire g6052;
wire II40594;
wire g28945;
wire g11590;
wire g16489;
wire g24140;
wire g25371;
wire g30751;
wire g29766;
wire g30945;
wire g8536;
wire g29980;
wire g9763;
wire g10460;
wire II17822;
wire g24834;
wire II40224;
wire g24940;
wire II24407;
wire g16505;
wire II39948;
wire g28315;
wire g16428;
wire g30117;
wire g13957;
wire II22679;
wire II14006;
wire g10810;
wire g5799;
wire g23846;
wire g11713;
wire g13221;
wire II33897;
wire II23380;
wire II14562;
wire g19664;
wire g21303;
wire II21083;
wire gbuf34;
wire II17801;
wire g27462;
wire g24821;
wire g21505;
wire II21389;
wire g28326;
wire g29488;
wire g16474;
wire g24442;
wire g24285;
wire g23066;
wire g11597;
wire II40760;
wire g11101;
wire g18505;
wire II24179;
wire II30810;
wire g23851;
wire g29434;
wire g15726;
wire II27346;
wire g28262;
wire II19605;
wire g16590;
wire g27034;
wire g18970;
wire II28813;
wire g28426;
wire g21800;
wire g14090;
wire g29378;
wire II28518;
wire g19839;
wire g8013;
wire g6289;
wire g28731;
wire g22126;
wire g9908;
wire g23167;
wire g21024;
wire g25830;
wire g21204;
wire g25064;
wire g9931;
wire g23177;
wire g25763;
wire II16153;
wire g25853;
wire g25444;
wire II29727;
wire g11948;
wire II18175;
wire g20402;
wire II20351;
wire g24312;
wire II21844;
wire gbuf213;
wire g26757;
wire g9664;
wire II40155;
wire g18718;
wire II14182;
wire g19052;
wire g5980;
wire II31781;
wire g19243;
wire g26167;
wire g13169;
wire g23241;
wire gbuf120;
wire g19067;
wire g13581;
wire g10113;
wire g6059;
wire g27936;
wire gbuf181;
wire II16300;
wire g18728;
wire g19692;
wire II30544;
wire g15508;
wire g10205;
wire g12349;
wire g28035;
wire g11078;
wire g17896;
wire g21253;
wire II16089;
wire g22634;
wire g11882;
wire g29517;
wire II24234;
wire II27260;
wire g12088;
wire g20431;
wire II23131;
wire g25295;
wire II25578;
wire II29415;
wire g27657;
wire II35905;
wire II23243;
wire II29625;
wire II23748;
wire II13190;
wire II18449;
wire g24506;
wire II25623;
wire g9760;
wire g17339;
wire g5754;
wire g30809;
wire g24164;
wire II13203;
wire g28072;
wire g26750;
wire g15128;
wire II34146;
wire II22572;
wire g19824;
wire g10555;
wire g24145;
wire g27142;
wire g24473;
wire II14547;
wire II29542;
wire II32943;
wire II13417;
wire II36568;
wire II13197;
wire g18951;
wire g18984;
wire g20369;
wire II31580;
wire g28013;
wire g25987;
wire g13512;
wire g10368;
wire II19938;
wire g27528;
wire II14660;
wire II24443;
wire g29853;
wire II23055;
wire g24553;
wire g5034;
wire g16322;
wire g22206;
wire g10283;
wire g15355;
wire g4498;
wire g11348;
wire II19645;
wire g25102;
wire II18106;
wire II26112;
wire II23226;
wire g10109;
wire g30641;
wire g11042;
wire g28414;
wire g26380;
wire g4794;
wire g8637;
wire g4191;
wire g19416;
wire g30648;
wire g30282;
wire g11555;
wire g24922;
wire g10161;
wire II34150;
wire gbuf85;
wire g22870;
wire g30292;
wire g27339;
wire g27174;
wire II31862;
wire II17066;
wire g15020;
wire II18288;
wire g29169;
wire g10337;
wire g23106;
wire g25887;
wire II20483;
wire g19020;
wire II31886;
wire g23513;
wire II39332;
wire g24252;
wire g27232;
wire II30305;
wire g5598;
wire g26063;
wire g15628;
wire II18835;
wire g4691;
wire g19847;
wire II40865;
wire II24215;
wire g24532;
wire II15642;
wire II25426;
wire g15560;
wire g15306;
wire II15935;
wire II34833;
wire II16587;
wire g29668;
wire g14691;
wire g25429;
wire II21246;
wire g30843;
wire g5591;
wire II24028;
wire g14541;
wire II23335;
wire II34456;
wire g19285;
wire g12003;
wire II16601;
wire g27981;
wire II32560;
wire II24709;
wire g10643;
wire g7466;
wire II28080;
wire g20114;
wire II19800;
wire g13096;
wire gbuf61;
wire II14243;
wire g22838;
wire g13648;
wire g12420;
wire g25941;
wire g29027;
wire g11085;
wire II40140;
wire g21864;
wire g24159;
wire g19741;
wire g10070;
wire g17798;
wire II28765;
wire g26002;
wire g19008;
wire g12545;
wire g14071;
wire g24576;
wire II36545;
wire g18295;
wire g28689;
wire g26813;
wire II29827;
wire g9301;
wire II13155;
wire g30942;
wire g21155;
wire g18915;
wire g13331;
wire g24798;
wire g18959;
wire g28750;
wire g27332;
wire g26525;
wire II27161;
wire g12502;
wire g21763;
wire g10327;
wire g21241;
wire g9440;
wire g15760;
wire II18359;
wire g30693;
wire g22082;
wire g25998;
wire g26987;
wire g21230;
wire g5606;
wire II23162;
wire g16705;
wire g26353;
wire g22273;
wire g23036;
wire II23651;
wire g5927;
wire g8493;
wire g25620;
wire g29695;
wire g17183;
wire g12523;
wire g7013;
wire g16357;
wire gbuf147;
wire g10041;
wire g23213;
wire II32468;
wire g30531;
wire g14450;
wire g21917;
wire II37765;
wire g28170;
wire g13417;
wire g29132;
wire g28429;
wire g29140;
wire g23971;
wire g20109;
wire g24624;
wire g11367;
wire g13412;
wire II17960;
wire g23140;
wire II32540;
wire g4286;
wire g30203;
wire gbuf134;
wire g7782;
wire II16880;
wire II36138;
wire g15569;
wire II18282;
wire II36230;
wire g29643;
wire gbuf25;
wire g25210;
wire g30482;
wire g23395;
wire g30662;
wire g15324;
wire g13774;
wire g28375;
wire g20963;
wire g20409;
wire II24444;
wire g7335;
wire g30401;
wire II31907;
wire g26577;
wire g28366;
wire g3521;
wire g15671;
wire g5959;
wire g13222;
wire g17664;
wire g28794;
wire g30767;
wire II35254;
wire g10529;
wire g19821;
wire II21505;
wire II14402;
wire g20704;
wire g8330;
wire g29578;
wire g16857;
wire g26776;
wire II36008;
wire g16189;
wire g24606;
wire II31387;
wire II41135;
wire gbuf163;
wire g5162;
wire II38833;
wire g15432;
wire II26512;
wire g15003;
wire g23271;
wire g5410;
wire g5817;
wire II31733;
wire g29615;
wire g25948;
wire II39863;
wire II20598;
wire g16105;
wire g23736;
wire II21918;
wire g9365;
wire g20769;
wire g24746;
wire g17924;
wire g20471;
wire g8339;
wire g11983;
wire g12850;
wire g14684;
wire g22174;
wire g22798;
wire g29204;
wire II41132;
wire g23162;
wire g14592;
wire g30065;
wire II23648;
wire II38860;
wire g22809;
wire II38125;
wire g9639;
wire g30744;
wire g10213;
wire g20449;
wire g9187;
wire g24876;
wire II39053;
wire g15282;
wire g22047;
wire g23136;
wire g16371;
wire II35852;
wire g29162;
wire II24537;
wire g29248;
wire g22627;
wire g22099;
wire g23568;
wire II32170;
wire II29802;
wire g9173;
wire II18432;
wire g19725;
wire g7548;
wire g22421;
wire g16761;
wire II40703;
wire g23979;
wire g26552;
wire g28674;
wire II38380;
wire g22755;
wire II15680;
wire g5826;
wire g28003;
wire g12747;
wire g27791;
wire II18464;
wire g19655;
wire g19454;
wire II18605;
wire II18438;
wire g9501;
wire g29074;
wire g9443;
wire II33570;
wire g25536;
wire g20900;
wire g10846;
wire g23137;
wire g17736;
wire II18160;
wire g26876;
wire II32642;
wire g13424;
wire g22997;
wire g29901;
wire g25074;
wire g15474;
wire II29259;
wire g25094;
wire g16878;
wire II35116;
wire g24613;
wire g6134;
wire g7639;
wire g15499;
wire g10168;
wire II40904;
wire g13027;
wire g5249;
wire II14040;
wire g7561;
wire g4913;
wire g19283;
wire g14131;
wire II36848;
wire II38838;
wire g29277;
wire g28149;
wire II33676;
wire g24358;
wire g5732;
wire II14755;
wire g16432;
wire g11874;
wire g13902;
wire g30441;
wire II37934;
wire g4520;
wire g10046;
wire g20882;
wire II40991;
wire g5402;
wire g30133;
wire g18265;
wire g28978;
wire g21284;
wire II19345;
wire II33586;
wire II25778;
wire g23885;
wire g8519;
wire g19629;
wire g11812;
wire g30224;
wire g29634;
wire g28889;
wire g26739;
wire g11505;
wire II29280;
wire g26010;
wire II20535;
wire g24343;
wire g5985;
wire g19740;
wire g3934;
wire g29665;
wire g27617;
wire g8494;
wire g29614;
wire g8387;
wire II39423;
wire g12554;
wire g22717;
wire g21610;
wire g28841;
wire g4936;
wire g9580;
wire II40269;
wire g19087;
wire g28711;
wire II14280;
wire g28659;
wire g4251;
wire II29345;
wire g27428;
wire II35470;
wire II29421;
wire g14268;
wire g30824;
wire II23698;
wire g4780;
wire g30106;
wire g18404;
wire g22730;
wire g26659;
wire g28849;
wire g19221;
wire g30388;
wire II31136;
wire g23075;
wire g11765;
wire g28165;
wire g27073;
wire g25118;
wire II30053;
wire g29572;
wire g18502;
wire g19043;
wire g19724;
wire g4982;
wire II36084;
wire II36256;
wire II36708;
wire g26496;
wire g12070;
wire g27872;
wire g16032;
wire II29933;
wire g26858;
wire g25805;
wire g28033;
wire g20926;
wire gbuf174;
wire II24521;
wire g19849;
wire g30721;
wire g29178;
wire g25658;
wire g27334;
wire g22067;
wire g22318;
wire g22261;
wire II30155;
wire g11321;
wire g10703;
wire II37185;
wire II25802;
wire II14742;
wire g22518;
wire g10706;
wire g13193;
wire II37050;
wire g21441;
wire g9724;
wire g3897;
wire g26713;
wire g15018;
wire II32844;
wire g10208;
wire g5115;
wire g22175;
wire g28066;
wire g21319;
wire II31577;
wire II24501;
wire g26703;
wire g23560;
wire g21749;
wire g19818;
wire g15143;
wire II36912;
wire II39985;
wire g15510;
wire g22265;
wire II23341;
wire g17271;
wire g30094;
wire g12960;
wire II35930;
wire II28825;
wire g21796;
wire g22229;
wire g8504;
wire g8183;
wire II26868;
wire g25250;
wire g23559;
wire g21314;
wire II34153;
wire II32874;
wire g8088;
wire g28779;
wire g27292;
wire II36150;
wire g30471;
wire g24745;
wire II35042;
wire g11533;
wire g28440;
wire g13145;
wire g17636;
wire g30325;
wire g24901;
wire g19762;
wire II33293;
wire g30023;
wire II21520;
wire g4475;
wire II33876;
wire II40481;
wire g18025;
wire II23754;
wire g11831;
wire g24430;
wire g13429;
wire g22249;
wire II35494;
wire g22341;
wire g5918;
wire II14529;
wire g30760;
wire g19634;
wire g24181;
wire g14985;
wire g18743;
wire II20553;
wire II38166;
wire g30097;
wire II28628;
wire g12807;
wire II16453;
wire II38936;
wire g20186;
wire g8551;
wire II17863;
wire g27732;
wire g18990;
wire II36105;
wire II23234;
wire g21310;
wire II29724;
wire g20464;
wire g7958;
wire g22224;
wire II31895;
wire g30270;
wire g21250;
wire g28675;
wire g21557;
wire g18892;
wire g5810;
wire g11151;
wire g23998;
wire II21959;
wire g12154;
wire g27432;
wire g19317;
wire g13557;
wire g30625;
wire g24720;
wire g27459;
wire II24178;
wire g22906;
wire g23235;
wire II21318;
wire g26732;
wire II35301;
wire g17270;
wire g26636;
wire II32854;
wire g23997;
wire g21799;
wire g10235;
wire g25619;
wire g29935;
wire g10077;
wire g23455;
wire g20246;
wire g12926;
wire II39782;
wire g18691;
wire g19558;
wire g19148;
wire g21063;
wire g20611;
wire g5932;
wire g26362;
wire g25122;
wire g21792;
wire g10407;
wire g13865;
wire g24373;
wire g20281;
wire II35124;
wire g22962;
wire g15774;
wire II30860;
wire II21407;
wire g16350;
wire g24854;
wire II29697;
wire II40131;
wire II18226;
wire g11749;
wire II20347;
wire g13186;
wire g29679;
wire g7876;
wire g28101;
wire g24941;
wire II32153;
wire g16894;
wire g12307;
wire g4962;
wire g24663;
wire g12048;
wire g24711;
wire II16044;
wire II31919;
wire g5876;
wire II37038;
wire II36240;
wire g22655;
wire g7872;
wire g19840;
wire g21952;
wire g29050;
wire g9026;
wire g10095;
wire g29241;
wire g23670;
wire II30925;
wire g22692;
wire II37083;
wire II25750;
wire g29345;
wire II27672;
wire g16993;
wire g27785;
wire II25474;
wire II24530;
wire g30155;
wire g23055;
wire g17936;
wire g11444;
wire II40294;
wire g25554;
wire g22289;
wire II32569;
wire II15222;
wire II35521;
wire g26674;
wire g17463;
wire g5893;
wire g25220;
wire g19153;
wire II39797;
wire II38378;
wire g13070;
wire g17132;
wire II23821;
wire II26940;
wire g27736;
wire g20793;
wire g8707;
wire g27956;
wire g24569;
wire II39776;
wire g8879;
wire II28564;
wire g18195;
wire g13941;
wire g4828;
wire g26616;
wire g20632;
wire g16493;
wire II25829;
wire g29101;
wire II31676;
wire g30035;
wire g20827;
wire g21129;
wire g25286;
wire g27134;
wire g9912;
wire g30511;
wire g8813;
wire II25921;
wire II22512;
wire g23621;
wire g16840;
wire II27107;
wire g28582;
wire g29553;
wire II39168;
wire g25865;
wire g29680;
wire II35961;
wire g26953;
wire II34791;
wire g22480;
wire g29100;
wire g13232;
wire g11905;
wire g21044;
wire g16201;
wire g28058;
wire g25634;
wire g10218;
wire g12942;
wire g15244;
wire g23317;
wire g27568;
wire g30555;
wire g21523;
wire g13386;
wire II29672;
wire II38878;
wire g23079;
wire g21926;
wire g562;
wire g22941;
wire g25343;
wire g9898;
wire g22748;
wire II16873;
wire II28090;
wire II35689;
wire g21167;
wire g29916;
wire II36894;
wire g8840;
wire g13870;
wire g12332;
wire II40970;
wire g7967;
wire g21095;
wire g25646;
wire g30708;
wire g13212;
wire g22338;
wire g10477;
wire g23905;
wire II40078;
wire g19225;
wire II17698;
wire g24695;
wire g13673;
wire g11894;
wire g30306;
wire g23501;
wire g27724;
wire g12768;
wire II38602;
wire II20625;
wire II30122;
wire II32607;
wire II36604;
wire g11868;
wire II16082;
wire II31460;
wire g29209;
wire II28034;
wire g7579;
wire g11779;
wire g20922;
wire II29174;
wire II19432;
wire g12105;
wire II27206;
wire g10127;
wire g27011;
wire g15476;
wire g22477;
wire g10293;
wire g26513;
wire g26433;
wire g23680;
wire II24485;
wire g13173;
wire g23598;
wire g18666;
wire g5092;
wire g11771;
wire g30735;
wire II18749;
wire II28305;
wire g27327;
wire II34476;
wire g22953;
wire g26272;
wire g16136;
wire g15834;
wire g8822;
wire g20355;
wire II27361;
wire g29799;
wire g25566;
wire g28356;
wire g26799;
wire g28229;
wire g13068;
wire g5352;
wire II35944;
wire g18861;
wire g23662;
wire g4130;
wire g25540;
wire g21711;
wire g23099;
wire g28456;
wire g16342;
wire g28647;
wire II22533;
wire II13095;
wire II31520;
wire g29534;
wire g8321;
wire g27216;
wire II26078;
wire II35503;
wire II24037;
wire g27448;
wire g6163;
wire II18052;
wire g17381;
wire g10615;
wire g11354;
wire g17913;
wire g30355;
wire II36574;
wire II25141;
wire g11432;
wire g27042;
wire g13637;
wire g19121;
wire g19703;
wire g10826;
wire g13310;
wire II19921;
wire g24867;
wire g20746;
wire g27146;
wire II14073;
wire g28083;
wire g23839;
wire II25847;
wire g26289;
wire g25039;
wire II31065;
wire g29549;
wire g19000;
wire g28155;
wire g11724;
wire g26341;
wire g10016;
wire g27358;
wire g13279;
wire g26956;
wire g22296;
wire g13309;
wire g20435;
wire g9401;
wire g28854;
wire II26654;
wire g12912;
wire g4375;
wire g16457;
wire g12159;
wire g23202;
wire II40733;
wire g29062;
wire II38689;
wire g29366;
wire g13043;
wire g18124;
wire g8472;
wire II27827;
wire II37784;
wire II40835;
wire II21647;
wire g24129;
wire g10220;
wire II35695;
wire g29272;
wire g27585;
wire g24453;
wire g9446;
wire g12418;
wire II30976;
wire II14877;
wire g30260;
wire II25303;
wire II27113;
wire g9094;
wire g16728;
wire g22770;
wire II25030;
wire g21699;
wire II14014;
wire g23689;
wire g18878;
wire II37593;
wire g8179;
wire g13105;
wire g30861;
wire g30312;
wire II19654;
wire g11547;
wire g16954;
wire g20118;
wire II18680;
wire g24126;
wire g23741;
wire g18038;
wire g24464;
wire g28387;
wire g30703;
wire gbuf98;
wire II30701;
wire II27324;
wire g20105;
wire g30000;
wire g23045;
wire g12050;
wire g5897;
wire g12275;
wire g11066;
wire II25810;
wire g11897;
wire g19531;
wire g18943;
wire g21461;
wire g27287;
wire g16853;
wire g16041;
wire g13465;
wire g10436;
wire II16900;
wire II26464;
wire g30015;
wire II35437;
wire II24655;
wire II27772;
wire g26189;
wire g8847;
wire g23936;
wire g24301;
wire II32577;
wire II30083;
wire II14984;
wire g15437;
wire II24513;
wire g27410;
wire g22743;
wire g26584;
wire g24101;
wire gbuf14;
wire II24381;
wire g12057;
wire g19511;
wire II30074;
wire g26921;
wire g25438;
wire II25633;
wire g26599;
wire g24593;
wire g23262;
wire g29413;
wire g8993;
wire II40814;
wire II39151;
wire g12447;
wire g15486;
wire g15376;
wire g22702;
wire g8910;
wire g21048;
wire g19180;
wire II22626;
wire g29694;
wire g29375;
wire g15931;
wire g10419;
wire II32184;
wire II16074;
wire g18275;
wire II24388;
wire g11841;
wire II38635;
wire g28345;
wire g8632;
wire g30800;
wire g9138;
wire II39017;
wire II23448;
wire g11166;
wire g23204;
wire g13894;
wire g26911;
wire II30179;
wire g20383;
wire g17360;
wire g17450;
wire II14799;
wire II23463;
wire II37041;
wire g24793;
wire g21292;
wire g18882;
wire g23070;
wire g12064;
wire g12150;
wire II20873;
wire g13624;
wire g15992;
wire g28963;
wire II20697;
wire g22846;
wire g27056;
wire g28758;
wire II34198;
wire g17830;
wire g29094;
wire g12969;
wire g10074;
wire II38011;
wire g29418;
wire II15899;
wire g19478;
wire g5646;
wire g3987;
wire g25772;
wire II33154;
wire g19754;
wire g18324;
wire g19882;
wire g18871;
wire II25108;
wire II39532;
wire g9082;
wire g21378;
wire II32634;
wire g26114;
wire g23209;
wire g8391;
wire g15573;
wire g24810;
wire II37982;
wire g16285;
wire g19671;
wire g13669;
wire II18031;
wire II30296;
wire g9484;
wire II33732;
wire g27149;
wire g23583;
wire g27163;
wire II38046;
wire g28447;
wire g26642;
wire g24235;
wire g14736;
wire g27371;
wire g17330;
wire II22962;
wire g26983;
wire II18728;
wire g24213;
wire g30697;
wire g5901;
wire g12302;
wire g21235;
wire g30561;
wire g14584;
wire g5710;
wire II30314;
wire g5871;
wire g28763;
wire g28724;
wire g24382;
wire g11968;
wire g25335;
wire g19165;
wire g6290;
wire g24723;
wire g29009;
wire g24774;
wire g14086;
wire g24336;
wire g29358;
wire g18834;
wire g28061;
wire g5556;
wire II37191;
wire g5764;
wire g12210;
wire g10196;
wire g22169;
wire II35868;
wire g20633;
wire g13141;
wire g19100;
wire g18765;
wire g7623;
wire II32724;
wire g25868;
wire g24109;
wire g20596;
wire g10171;
wire g5920;
wire II29575;
wire g28252;
wire g30217;
wire g27553;
wire II23567;
wire g27534;
wire g23798;
wire II18701;
wire g19150;
wire II40667;
wire II40320;
wire g23082;
wire g20607;
wire g18587;
wire II15958;
wire II23968;
wire II35772;
wire g24514;
wire g23187;
wire g6098;
wire g12263;
wire g30163;
wire II30568;
wire II19485;
wire II29975;
wire g23186;
wire g29786;
wire g12487;
wire II25129;
wire g28008;
wire g26434;
wire II15978;
wire II40179;
wire g22831;
wire g26885;
wire g21660;
wire II26596;
wire g20314;
wire g17599;
wire g19174;
wire II21286;
wire g24817;
wire g25338;
wire g13130;
wire g27824;
wire II35919;
wire g29877;
wire II28229;
wire II24394;
wire II23074;
wire II24626;
wire g4651;
wire II28051;
wire g28094;
wire gbuf201;
wire II25732;
wire II27212;
wire g8221;
wire g26532;
wire g10476;
wire g9383;
wire II38695;
wire g20468;
wire g10444;
wire g6027;
wire g21016;
wire g18989;
wire g30070;
wire g26600;
wire g20612;
wire g4641;
wire g10804;
wire g18606;
wire g20459;
wire II40889;
wire g20903;
wire g21021;
wire g22217;
wire g28105;
wire II24913;
wire g9759;
wire II17966;
wire g19060;
wire gbuf91;
wire II17872;
wire gbuf52;
wire g21959;
wire II22828;
wire g11376;
wire g30921;
wire g10371;
wire g5409;
wire II31628;
wire g19921;
wire II24194;
wire g20640;
wire II16150;
wire g22074;
wire g8440;
wire g28783;
wire g27047;
wire g20148;
wire II25721;
wire g4544;
wire g20875;
wire II31688;
wire g4647;
wire II39622;
wire g27667;
wire g17506;
wire II33867;
wire g21995;
wire g9462;
wire g6180;
wire g17222;
wire g27718;
wire g28321;
wire g16616;
wire g21270;
wire g14718;
wire II31601;
wire g10465;
wire g23605;
wire II30552;
wire II39404;
wire g21361;
wire g8554;
wire g19334;
wire g8545;
wire g8098;
wire g23633;
wire g24418;
wire g9248;
wire g22824;
wire g9479;
wire g26663;
wire g5543;
wire II37725;
wire II36676;
wire II32102;
wire g28391;
wire g15820;
wire g9756;
wire gbuf208;
wire g10461;
wire g5255;
wire II23451;
wire g24826;
wire g14366;
wire g8835;
wire gbuf177;
wire g22640;
wire g27120;
wire g11991;
wire g10118;
wire g17543;
wire II34659;
wire II24076;
wire II19702;
wire II36738;
wire g22202;
wire g17057;
wire g30928;
wire g27230;
wire g30540;
wire g25133;
wire g30267;
wire g28709;
wire g22623;
wire II38641;
wire II31904;
wire II33421;
wire g21842;
wire g25368;
wire II37324;
wire g17903;
wire g21457;
wire g22789;
wire g30470;
wire II23958;
wire g30656;
wire g22408;
wire g10048;
wire g22367;
wire g30079;
wire g28540;
wire II37176;
wire g25402;
wire g29156;
wire II31589;
wire g19041;
wire g21700;
wire g16515;
wire II40071;
wire g24962;
wire g13449;
wire g27768;
wire g30456;
wire g17887;
wire g28398;
wire g13882;
wire g18863;
wire g17601;
wire II38975;
wire II28133;
wire g20127;
wire g30126;
wire g5272;
wire g24110;
wire g12231;
wire g11465;
wire g4098;
wire g22034;
wire g22240;
wire II35890;
wire g23866;
wire g22015;
wire g28431;
wire g21786;
wire g18962;
wire II20959;
wire g27095;
wire g30299;
wire g30570;
wire g19113;
wire g9505;
wire g19480;
wire g26542;
wire g18877;
wire II40170;
wire g10995;
wire II23105;
wire g6887;
wire II17978;
wire g11863;
wire g26191;
wire II23253;
wire g13858;
wire g5998;
wire II22974;
wire II14811;
wire II13907;
wire II17677;
wire II39899;
wire g21778;
wire g7970;
wire g21393;
wire g29525;
wire g10595;
wire II21769;
wire g25030;
wire g30468;
wire g22886;
wire g29648;
wire gbuf159;
wire II18399;
wire g25838;
wire g8894;
wire II36673;
wire g12076;
wire II22768;
wire II15964;
wire g6638;
wire g5978;
wire g24066;
wire g15336;
wire g20555;
wire II29087;
wire g19214;
wire g23304;
wire g29453;
wire II16292;
wire g15524;
wire g20013;
wire g18831;
wire g19813;
wire g30538;
wire g27254;
wire g15801;
wire g30515;
wire II13919;
wire II39843;
wire g23192;
wire II34204;
wire g11816;
wire g20979;
wire g19385;
wire g12995;
wire II17666;
wire II29957;
wire II30838;
wire g23193;
wire II36300;
wire g22304;
wire g12923;
wire g21473;
wire g22021;
wire g13158;
wire g10184;
wire g13242;
wire g19755;
wire g22734;
wire g24349;
wire g26216;
wire g25880;
wire g16692;
wire g18312;
wire g29312;
wire g22763;
wire g28339;
wire g11976;
wire g28651;
wire II30044;
wire g30981;
wire II26567;
wire II25300;
wire II14037;
wire g20325;
wire g10313;
wire g29083;
wire g21194;
wire g26791;
wire II24102;
wire g16449;
wire g26787;
wire g27889;
wire g9101;
wire g24447;
wire gbuf37;
wire g10509;
wire g21418;
wire g15349;
wire g22497;
wire g29991;
wire g26358;
wire g25675;
wire g10266;
wire g9439;
wire II33695;
wire II35017;
wire g22713;
wire g23619;
wire g6061;
wire g19388;
wire g10249;
wire g21960;
wire g26607;
wire g22792;
wire II25534;
wire g22723;
wire g9923;
wire g30398;
wire g24803;
wire II32716;
wire g5885;
wire II38707;
wire II20655;
wire g20254;
wire g17227;
wire II24416;
wire g11636;
wire II16009;
wire II41019;
wire II39812;
wire g6037;
wire II28455;
wire g29551;
wire g15142;
wire g29160;
wire g20395;
wire g12017;
wire g28378;
wire II33589;
wire g10257;
wire g3948;
wire g24477;
wire g8853;
wire g20444;
wire g25346;
wire g28491;
wire g30954;
wire g30259;
wire II25516;
wire g29238;
wire II23161;
wire II25291;
wire g3245;
wire g29801;
wire II18022;
wire II16347;
wire g25091;
wire g29341;
wire g23829;
wire II37846;
wire g13560;
wire g8411;
wire g13390;
wire g28551;
wire II40263;
wire II32587;
wire g17197;
wire II25701;
wire g21536;
wire g13269;
wire g24845;
wire II36978;
wire g28234;
wire g25229;
wire g28679;
wire g9196;
wire g25166;
wire gbuf170;
wire g10024;
wire II14937;
wire g9518;
wire g8805;
wire II18347;
wire g27539;
wire g19452;
wire g9145;
wire II23709;
wire g13215;
wire g24141;
wire g14052;
wire II35464;
wire g21681;
wire g26473;
wire g21322;
wire g12451;
wire g14273;
wire g16558;
wire g13341;
wire g16001;
wire g22040;
wire II21190;
wire g29423;
wire II18178;
wire II31661;
wire g12253;
wire g30362;
wire g6631;
wire g5861;
wire II18842;
wire g21054;
wire g29732;
wire II37023;
wire II35034;
wire II31436;
wire II35974;
wire g21398;
wire g5966;
wire II24695;
wire g24174;
wire g24761;
wire II31024;
wire g24797;
wire II29585;
wire II35482;
wire II17303;
wire II33726;
wire g12285;
wire g12139;
wire g12857;
wire g14022;
wire g8567;
wire g4392;
wire g13209;
wire g15461;
wire II31144;
wire II35859;
wire g9885;
wire II35422;
wire g7912;
wire II16283;
wire g29969;
wire g19606;
wire g10151;
wire g16501;
wire g9066;
wire g23548;
wire g25329;
wire II21127;
wire II19718;
wire g8751;
wire g5647;
wire II30158;
wire g9498;
wire g21112;
wire II22521;
wire g11805;
wire g20372;
wire g29252;
wire g25787;
wire g25154;
wire II35976;
wire g13488;
wire g13115;
wire g4176;
wire g27242;
wire g16184;
wire g29951;
wire g24130;
wire g21368;
wire g19145;
wire g11173;
wire g27195;
wire g17174;
wire g13538;
wire II40790;
wire II18722;
wire g17076;
wire g24329;
wire II37284;
wire II22800;
wire g15730;
wire g17430;
wire g10381;
wire g9004;
wire g26694;
wire g15049;
wire g16498;
wire II22885;
wire II22803;
wire g4581;
wire g30408;
wire g28650;
wire g3566;
wire II35993;
wire g6676;
wire g24221;
wire g6418;
wire g16098;
wire g26546;
wire II31502;
wire g10891;
wire g27382;
wire II27281;
wire g26678;
wire g11718;
wire II17780;
wire g22865;
wire II36592;
wire g22257;
wire II33327;
wire g13481;
wire g25219;
wire II32462;
wire g16764;
wire g26561;
wire g20305;
wire g22337;
wire II40847;
wire g10004;
wire g30274;
wire II19971;
wire II22506;
wire g7652;
wire g25264;
wire g11823;
wire g4787;
wire g4602;
wire g10067;
wire g10773;
wire g19303;
wire g28493;
wire g17262;
wire g12608;
wire II21803;
wire II37303;
wire g10532;
wire g28188;
wire g16302;
wire II39273;
wire g21759;
wire g12117;
wire g5361;
wire II27379;
wire II36301;
wire g16119;
wire g20943;
wire gbuf106;
wire g22659;
wire g15764;
wire g29558;
wire g11420;
wire g9770;
wire II37991;
wire g19448;
wire g20377;
wire g19037;
wire II38196;
wire g6209;
wire g22253;
wire g19234;
wire g25847;
wire g13868;
wire g13325;
wire g29509;
wire g23740;
wire II38071;
wire g15139;
wire II37029;
wire g21382;
wire II37566;
wire II40039;
wire g25928;
wire g20484;
wire g18485;
wire II34993;
wire II23608;
wire g14966;
wire g10677;
wire g13500;
wire g28308;
wire II17998;
wire g30883;
wire g5926;
wire g7919;
wire g22197;
wire g18848;
wire g16864;
wire g18944;
wire g9110;
wire g22056;
wire II36744;
wire g25798;
wire g17448;
wire g4234;
wire g14292;
wire II32964;
wire g16055;
wire g7471;
wire II33711;
wire g21553;
wire g18110;
wire g26372;
wire g23918;
wire g23147;
wire g24273;
wire II21449;
wire II29339;
wire g16368;
wire g10057;
wire g17788;
wire g5868;
wire g22523;
wire g27329;
wire II27917;
wire g20458;
wire II41012;
wire g21902;
wire g11091;
wire g11797;
wire g27704;
wire g30892;
wire II24531;
wire g23612;
wire g20286;
wire g18553;
wire II15613;
wire II15998;
wire g28095;
wire g29448;
wire II26051;
wire g9592;
wire g26314;
wire II20816;
wire g5809;
wire g22769;
wire II34674;
wire g12160;
wire g11959;
wire II18515;
wire g30498;
wire g7559;
wire g25417;
wire g18783;
wire g8465;
wire g21325;
wire II30864;
wire g6146;
wire gbuf160;
wire II36496;
wire g14577;
wire g27341;
wire g10946;
wire g29956;
wire II33804;
wire g30507;
wire g18824;
wire II16432;
wire g29949;
wire g11549;
wire II17875;
wire g15639;
wire g15902;
wire g28481;
wire g15582;
wire g12195;
wire II17746;
wire g26807;
wire g14954;
wire g26293;
wire g23144;
wire g22786;
wire g8548;
wire g28624;
wire g10673;
wire g11733;
wire g19055;
wire g21860;
wire g28219;
wire g24097;
wire g20417;
wire g4153;
wire g13020;
wire g18927;
wire g9356;
wire g26044;
wire II14609;
wire g27994;
wire g5636;
wire g30347;
wire II13107;
wire g18996;
wire II13940;
wire g9416;
wire g11653;
wire II34809;
wire g11740;
wire g26235;
wire g25324;
wire II19634;
wire g26782;
wire II40910;
wire g25238;
wire g15970;
wire g10120;
wire II20009;
wire II17795;
wire g30444;
wire g30321;
wire g4908;
wire g8103;
wire II15859;
wire II15212;
wire gbuf195;
wire g19099;
wire g23526;
wire g27574;
wire II15876;
wire II24015;
wire g29716;
wire g13135;
wire II16104;
wire g27300;
wire II31286;
wire II40501;
wire II39375;
wire g30855;
wire g29960;
wire g9016;
wire g27666;
wire g11228;
wire g30605;
wire g4529;
wire g26825;
wire g10693;
wire g19856;
wire g8696;
wire g10539;
wire g17714;
wire II30636;
wire II14760;
wire g29211;
wire g21714;
wire g13845;
wire g9780;
wire g17204;
wire g30084;
wire g22212;
wire II27275;
wire g10060;
wire g28749;
wire g19327;
wire II21974;
wire II32379;
wire g26015;
wire g6905;
wire II23067;
wire g27153;
wire II31547;
wire g18645;
wire II21612;
wire g13704;
wire g23635;
wire g5798;
wire II26437;
wire g28658;
wire g20608;
wire II37232;
wire g29180;
wire II30017;
wire g3998;
wire g29328;
wire II16967;
wire g11576;
wire g20772;
wire II14839;
wire g16129;
wire g24787;
wire g3975;
wire II20706;
wire g15574;
wire II33286;
wire g16849;
wire g10683;
wire II25938;
wire g27320;
wire g22180;
wire g11495;
wire g29635;
wire II25717;
wire II25791;
wire g4278;
wire g5665;
wire g8907;
wire II18127;
wire g21661;
wire g16966;
wire g24766;
wire g9170;
wire g17156;
wire g30411;
wire g16719;
wire g23723;
wire II15442;
wire g20390;
wire II32519;
wire g29106;
wire II25032;
wire II16444;
wire g30636;
wire g23463;
wire g18965;
wire g10086;
wire g22187;
wire g21943;
wire II36217;
wire II14602;
wire g17201;
wire g17853;
wire g6016;
wire g15789;
wire g29540;
wire II38360;
wire g22317;
wire II23180;
wire g4049;
wire II23103;
wire g29172;
wire II22937;
wire g4171;
wire g18140;
wire II23274;
wire II31946;
wire g26722;
wire g17814;
wire g12135;
wire g5707;
wire g8126;
wire g28403;
wire g26387;
wire g20492;
wire g19551;
wire II18262;
wire g18331;
wire g13992;
wire II16489;
wire g21726;
wire g9604;
wire g29088;
wire II32423;
wire g12012;
wire g19774;
wire g19320;
wire II15971;
wire g13181;
wire g28048;
wire g9648;
wire II34977;
wire g5296;
wire g27680;
wire g23886;
wire g21565;
wire g3925;
wire g26474;
wire II30119;
wire g30024;
wire II15204;
wire g9241;
wire II33643;
wire II41047;
wire g30489;
wire g23123;
wire g27108;
wire g22868;
wire II33708;
wire II20568;
wire g9810;
wire g10100;
wire g19588;
wire g27415;
wire g19567;
wire g30113;
wire g5702;
wire II20631;
wire II38480;
wire g23879;
wire g20786;
wire g3919;
wire g24308;
wire g11950;
wire g20197;
wire g29931;
wire g25615;
wire II23917;
wire II19791;
wire g27305;
wire II22509;
wire g27100;
wire g30977;
wire g12495;
wire g13438;
wire g23942;
wire II25389;
wire g23403;
wire g7533;
wire II23036;
wire g16005;
wire g17661;
wire g8515;
wire II35926;
wire g27367;
wire II29389;
wire II16002;
wire g11758;
wire g8481;
wire g4112;
wire g24562;
wire g20575;
wire g26033;
wire II36390;
wire g11937;
wire g23288;
wire g6119;
wire g15268;
wire g25045;
wire g24393;
wire II25653;
wire g25892;
wire g23006;
wire g28775;
wire g5961;
wire g15236;
wire g30813;
wire g29672;
wire g5413;
wire g24013;
wire g16028;
wire II23763;
wire g21389;
wire g16278;
wire II39011;
wire g19792;
wire g14201;
wire II25156;
wire g13198;
wire g4680;
wire g30056;
wire II15457;
wire g24933;
wire II23745;
wire II34746;
wire g14336;
wire g5942;
wire g30835;
wire g21814;
wire g8947;
wire II38599;
wire g25852;
wire g29811;
wire g21969;
wire II13965;
wire II17150;
wire II24555;
wire g10569;
wire II38755;
wire g30701;
wire II36921;
wire g12559;
wire II40239;
wire g22058;
wire g25172;
wire g20294;
wire g22333;
wire II16179;
wire g11862;
wire g21537;
wire g25436;
wire II33849;
wire II19689;
wire g26497;
wire g24127;
wire II31922;
wire g24354;
wire g14922;
wire II15398;
wire g13305;
wire II21064;
wire g22185;
wire g25191;
wire II30467;
wire g15172;
wire g4111;
wire II39457;
wire g8487;
wire II33703;
wire g16026;
wire g17410;
wire g19053;
wire g7555;
wire g15112;
wire II13211;
wire g15265;
wire g6034;
wire g21770;
wire g7570;
wire g23406;
wire II27059;
wire g7658;
wire II25914;
wire g28235;
wire II34743;
wire g25817;
wire g20531;
wire g24433;
wire g9621;
wire g13978;
wire g24248;
wire II30287;
wire g8278;
wire g8946;
wire g21967;
wire g29232;
wire g28112;
wire g27492;
wire g26728;
wire II30248;
wire II17632;
wire g10940;
wire II27080;
wire g23047;
wire g9338;
wire g28092;
wire II36984;
wire g26788;
wire II37605;
wire g19876;
wire g30476;
wire g18538;
wire g8084;
wire g25048;
wire g14337;
wire g27915;
wire g17812;
wire g26603;
wire g30532;
wire g20491;
wire g15231;
wire g23718;
wire g30458;
wire g26540;
wire g8801;
wire II38680;
wire g21090;
wire g21124;
wire g8468;
wire g10310;
wire g30772;
wire II37266;
wire g5778;
wire g5968;
wire g8904;
wire g9606;
wire g27301;
wire II23772;
wire II25186;
wire II27534;
wire g30791;
wire g23028;
wire II23154;
wire g9901;
wire gbuf10;
wire II14069;
wire II23545;
wire g18358;
wire g5283;
wire g28436;
wire g8941;
wire g30939;
wire II28346;
wire g28190;
wire g29103;
wire II38548;
wire g27809;
wire g4897;
wire II28984;
wire g9184;
wire g22178;
wire g23280;
wire g13113;
wire II16332;
wire g22063;
wire g16186;
wire II38363;
wire g22741;
wire g25873;
wire g13326;
wire g11259;
wire II21726;
wire g23468;
wire g24538;
wire g24059;
wire g29386;
wire g8717;
wire II30954;
wire g10877;
wire II18743;
wire II35702;
wire II19924;
wire g29542;
wire g6890;
wire g9809;
wire II36731;
wire g29921;
wire g25605;
wire II23418;
wire g11545;
wire II37116;
wire g10872;
wire II25386;
wire g27283;
wire g26684;
wire g15876;
wire g27530;
wire g16913;
wire g26646;
wire g3922;
wire g24340;
wire g30445;
wire II27089;
wire II36291;
wire II25889;
wire g27685;
wire II17866;
wire g26655;
wire II33840;
wire g12874;
wire II30489;
wire g4150;
wire g16910;
wire g20413;
wire g30328;
wire g9962;
wire g11980;
wire g10778;
wire g16387;
wire g26507;
wire II30227;
wire II36257;
wire g28836;
wire g26721;
wire g17055;
wire II36593;
wire II30170;
wire g11472;
wire g27800;
wire g20571;
wire g19631;
wire g30273;
wire II40826;
wire g13866;
wire g19868;
wire g16844;
wire II28369;
wire g21119;
wire g5318;
wire g22194;
wire g27107;
wire II23701;
wire g20822;
wire g14490;
wire g26091;
wire g16174;
wire II33906;
wire g15258;
wire g12116;
wire II40158;
wire g11818;
wire g18904;
wire g29145;
wire II20448;
wire g29710;
wire II34238;
wire g9665;
wire g28380;
wire II32109;
wire g15854;
wire g25126;
wire g29820;
wire g9276;
wire g12934;
wire g22756;
wire g24376;
wire gbuf89;
wire g28318;
wire g5135;
wire g15040;
wire g20880;
wire II40297;
wire g4899;
wire g29963;
wire g21327;
wire II19621;
wire g18786;
wire g22161;
wire II32042;
wire II34102;
wire g21928;
wire g12330;
wire II18533;
wire II36290;
wire g11575;
wire g13562;
wire g22971;
wire II31916;
wire II21939;
wire II26369;
wire g21072;
wire g27340;
wire II24104;
wire g25321;
wire g17839;
wire g4717;
wire g16850;
wire g24132;
wire II15288;
wire g28625;
wire g4127;
wire g19275;
wire g18257;
wire g17428;
wire g5947;
wire g29683;
wire g5946;
wire II30080;
wire g10125;
wire II39881;
wire II20744;
wire g14102;
wire g18925;
wire g11331;
wire g27939;
wire g6086;
wire g14642;
wire g11117;
wire g30845;
wire g29060;
wire g3990;
wire II16593;
wire g19858;
wire g11829;
wire g22903;
wire g12748;
wire g18164;
wire II16627;
wire II25728;
wire g28311;
wire g4925;
wire II32378;
wire II36078;
wire II16766;
wire g21944;
wire II18581;
wire g24594;
wire II32937;
wire g17753;
wire g29195;
wire g22966;
wire g14774;
wire g29349;
wire II32910;
wire g26656;
wire g27205;
wire g18993;
wire g16455;
wire g29652;
wire g27932;
wire g8044;
wire g18102;
wire g29938;
wire II15803;
wire g11284;
wire II31085;
wire II14449;
wire II27646;
wire g5512;
wire II30601;
wire g22122;
wire g21018;
wire g22031;
wire g28899;
wire g20537;
wire II13165;
wire g23039;
wire g25999;
wire II38758;
wire II40597;
wire g9868;
wire g21108;
wire g11954;
wire g27049;
wire II25595;
wire II38842;
wire g11032;
wire II15211;
wire g23061;
wire g25116;
wire II15556;
wire g13462;
wire g23909;
wire g24622;
wire g15412;
wire g19625;
wire II34313;
wire g26298;
wire II23725;
wire II38163;
wire g20917;
wire g26909;
wire g22356;
wire g20183;
wire g30316;
wire II20429;
wire g26626;
wire g16380;
wire g11633;
wire g12184;
wire II32518;
wire g19797;
wire II25862;
wire g23528;
wire II24577;
wire g26102;
wire g30558;
wire g12208;
wire g19544;
wire g9225;
wire II39065;
wire g11938;
wire g11953;
wire II30973;
wire II23833;
wire g17985;
wire g26401;
wire II31523;
wire g5906;
wire II24264;
wire g21530;
wire g10222;
wire g27093;
wire g22252;
wire g19590;
wire g10081;
wire II24017;
wire II13316;
wire II23279;
wire II32883;
wire II23510;
wire g15446;
wire g19934;
wire II27250;
wire g8227;
wire g12535;
wire g23659;
wire II33990;
wire II23655;
wire g17767;
wire g4249;
wire II34453;
wire g9374;
wire g24274;
wire II18151;
wire g20212;
wire g13484;
wire II13430;
wire g11613;
wire g23577;
wire gbuf82;
wire g20743;
wire II23018;
wire II24726;
wire g15352;
wire g24096;
wire g10527;
wire g8206;
wire g13505;
wire g20627;
wire g5820;
wire g13963;
wire g18847;
wire g21810;
wire g28208;
wire II29294;
wire g17181;
wire g10279;
wire g11163;
wire g4468;
wire g27244;
wire g5038;
wire g17967;
wire II16360;
wire g4508;
wire g28415;
wire g27193;
wire g16855;
wire g26034;
wire g18154;
wire II17278;
wire II23487;
wire g21178;
wire II31232;
wire g13271;
wire g30916;
wire g19306;
wire g24298;
wire II38202;
wire g21602;
wire g26520;
wire g30926;
wire II33460;
wire g15933;
wire II39533;
wire II31865;
wire II17557;
wire II14034;
wire II19750;
wire g17353;
wire g28207;
wire g10972;
wire g12643;
wire g7143;
wire II35313;
wire g13164;
wire g19216;
wire g11697;
wire g21148;
wire g11491;
wire g10152;
wire g25005;
wire II32150;
wire g21518;
wire g21741;
wire g22256;
wire II14532;
wire g26837;
wire g7593;
wire II37768;
wire II25249;
wire g20119;
wire II29073;
wire g23913;
wire g25017;
wire II38811;
wire g20588;
wire II31679;
wire II15863;
wire g10384;
wire g28682;
wire g22440;
wire g23772;
wire g13185;
wire g21304;
wire g16164;
wire g19503;
wire g20328;
wire II25207;
wire g29250;
wire II23507;
wire II17225;
wire g11820;
wire II14565;
wire g8891;
wire g23441;
wire g11764;
wire II23200;
wire g30602;
wire g4824;
wire g11931;
wire g19501;
wire g29941;
wire II18764;
wire g13210;
wire g18556;
wire g28496;
wire g10545;
wire g23676;
wire II34961;
wire g30628;
wire II40802;
wire g23724;
wire g19957;
wire g24384;
wire g29699;
wire g29805;
wire g30889;
wire g7461;
wire II25216;
wire g17534;
wire g20479;
wire II24765;
wire g25024;
wire g29342;
wire II24401;
wire II28450;
wire g16325;
wire g20051;
wire g28470;
wire g29739;
wire II13125;
wire g9876;
wire II18698;
wire g20394;
wire g8565;
wire g19918;
wire g26028;
wire g12136;
wire g17658;
wire g22867;
wire g28453;
wire g16093;
wire g12604;
wire g30110;
wire g27787;
wire g14955;
wire g29428;
wire g23259;
wire g12068;
wire g23113;
wire II30891;
wire g25196;
wire g26785;
wire g10692;
wire g5650;
wire II37790;
wire g20082;
wire g17225;
wire II17149;
wire g20102;
wire g19600;
wire g13202;
wire g22520;
wire g17876;
wire II20858;
wire II25021;
wire II23082;
wire II14641;
wire g30737;
wire g25244;
wire g5405;
wire g23856;
wire II17048;
wire g30706;
wire g5630;
wire II31850;
wire II25102;
wire g26993;
wire g4404;
wire g21707;
wire II32296;
wire g29554;
wire g17268;
wire g24652;
wire g26564;
wire g29444;
wire g17285;
wire II19503;
wire g30251;
wire g23545;
wire g26707;
wire g19776;
wire II41096;
wire II14094;
wire g26237;
wire g6064;
wire g21153;
wire g11857;
wire g10052;
wire g17815;
wire g16403;
wire g15136;
wire g4873;
wire g16567;
wire g21364;
wire II32710;
wire g29239;
wire g3945;
wire II18548;
wire g17588;
wire g11616;
wire II30209;
wire II30985;
wire g29022;
wire g25070;
wire g13507;
wire II22866;
wire g23824;
wire g22567;
wire g20707;
wire g24802;
wire II27270;
wire g14596;
wire g17030;
wire g8446;
wire II26843;
wire g25213;
wire g29188;
wire g9404;
wire g21495;
wire g18572;
wire g15408;
wire g29664;
wire g13430;
wire g4048;
wire g27879;
wire g21395;
wire g30750;
wire g29318;
wire g23613;
wire g25268;
wire g5882;
wire II31021;
wire g13003;
wire g5712;
wire II29098;
wire g11869;
wire II29101;
wire g21277;
wire g21766;
wire II17689;
wire g5138;
wire g11114;
wire g23779;
wire II21178;
wire g16560;
wire II23406;
wire g8501;
wire g14044;
wire g22794;
wire g19039;
wire g18840;
wire g21981;
wire II30611;
wire g19569;
wire g25301;
wire II33974;
wire II40952;
wire II23996;
wire g29773;
wire g29567;
wire g23615;
wire II22548;
wire g18593;
wire g24404;
wire g25169;
wire II29472;
wire g5864;
wire g18131;
wire g28330;
wire g29166;
wire g27708;
wire g16968;
wire g8540;
wire g16697;
wire g29451;
wire g5395;
wire g12909;
wire II17901;
wire II24327;
wire g5689;
wire g17640;
wire g25188;
wire II24669;
wire g28257;
wire g17474;
wire g28664;
wire g13983;
wire II29852;
wire g20939;
wire g27198;
wire g12992;
wire g25043;
wire g10977;
wire g29108;
wire g28328;
wire g24978;
wire g23865;
wire g29673;
wire g14032;
wire II28314;
wire g11358;
wire g20569;
wire g19814;
wire II33995;
wire g14668;
wire II37053;
wire g12449;
wire g30272;
wire II14769;
wire g11586;
wire g30789;
wire g23877;
wire g19176;
wire g26389;
wire g28260;
wire II40559;
wire gbuf108;
wire g11716;
wire g18967;
wire g28802;
wire g4044;
wire g5984;
wire g20131;
wire II35681;
wire g27713;
wire g27117;
wire g12086;
wire g4574;
wire g14256;
wire g19926;
wire II16141;
wire g23194;
wire g9124;
wire II21790;
wire II35434;
wire II18820;
wire g28683;
wire g18972;
wire g21848;
wire gbuf72;
wire g24683;
wire g23424;
wire g23349;
wire g11660;
wire g9595;
wire g7603;
wire g7482;
wire II14816;
wire II37623;
wire II30560;
wire II28096;
wire g25376;
wire g24216;
wire II27343;
wire II31604;
wire g15460;
wire g24231;
wire g23889;
wire g27659;
wire g13885;
wire g18879;
wire g19954;
wire g19709;
wire g29213;
wire g16665;
wire g18400;
wire g5693;
wire II23564;
wire II40964;
wire g11992;
wire II25625;
wire g30731;
wire g27725;
wire II29064;
wire g7972;
wire II37823;
wire g19236;
wire II34195;
wire g23686;
wire g17190;
wire g29135;
wire g19586;
wire gbuf183;
wire II19847;
wire g24458;
wire g9095;
wire II22022;
wire II31550;
wire II18046;
wire g8418;
wire g20558;
wire g28881;
wire g18809;
wire g13102;
wire II27395;
wire II24611;
wire g10440;
wire g4343;
wire g10507;
wire g28595;
wire II17238;
wire g18981;
wire g20553;
wire g19784;
wire g24167;
wire g5875;
wire g18236;
wire II32393;
wire II30290;
wire g10194;
wire g10536;
wire g21349;
wire g3833;
wire g12169;
wire g19047;
wire g29269;
wire g13945;
wire gbuf155;
wire g11557;
wire g7227;
wire gbuf171;
wire g20006;
wire g29526;
wire II22590;
wire g30356;
wire g11844;
wire g30076;
wire g24759;
wire g17620;
wire II38719;
wire g17545;
wire g27952;
wire g11306;
wire g28697;
wire g16068;
wire II31466;
wire g8846;
wire g9786;
wire g5547;
wire g23385;
wire II18010;
wire g21777;
wire g5087;
wire II32958;
wire g13109;
wire g24869;
wire II16608;
wire g26963;
wire g15105;
wire II31068;
wire g18521;
wire II33358;
wire g27258;
wire g15531;
wire g28012;
wire g16470;
wire g25330;
wire II27104;
wire g25290;
wire g22773;
wire II18752;
wire II15818;
wire g15819;
wire g11960;
wire II23954;
wire g13954;
wire g7531;
wire g25337;
wire g22873;
wire g16974;
wire II18172;
wire g8788;
wire g10624;
wire g16237;
wire g30718;
wire g19240;
wire II16241;
wire g11630;
wire II32470;
wire g12080;
wire g5346;
wire g25034;
wire g24814;
wire g23597;
wire g4650;
wire g13605;
wire g8681;
wire g13073;
wire II30841;
wire II36732;
wire g23217;
wire II29107;
wire II23739;
wire g30684;
wire g27092;
wire g8557;
wire II24092;
wire g21259;
wire g30840;
wire g21956;
wire II39252;
wire II23785;
wire g30366;
wire g4179;
wire g15771;
wire g20617;
wire II31646;
wire g5217;
wire g13861;
wire g18129;
wire g27780;
wire II30663;
wire g4601;
wire g6200;
wire g27009;
wire g26629;
wire g16639;
wire II40654;
wire gbuf30;
wire g10594;
wire g30103;
wire II14874;
wire II17122;
wire g26312;
wire g27347;
wire g15848;
wire g20381;
wire g15790;
wire g13240;
wire II27969;
wire g18891;
wire g19218;
wire g18548;
wire g12103;
wire g26183;
wire g27212;
wire g16250;
wire II16954;
wire g12920;
wire g26455;
wire II31658;
wire II17097;
wire g27126;
wire g22942;
wire g24780;
wire g4221;
wire II24226;
wire II32979;
wire g22278;
wire II39856;
wire g30286;
wire g10581;
wire II40757;
wire g28850;
wire g13847;
wire g24811;
wire g25137;
wire g22766;
wire g22133;
wire g26211;
wire g28722;
wire II18713;
wire g9956;
wire II36533;
wire g23307;
wire g10438;
wire II31682;
wire g22292;
wire g11723;
wire g25835;
wire g26846;
wire g19198;
wire g5995;
wire II17995;
wire g30147;
wire II21292;
wire II38401;
wire g29293;
wire II30854;
wire II20691;
wire g7157;
wire g30618;
wire g8550;
wire g14067;
wire II30089;
wire g14413;
wire II36316;
wire g20190;
wire g10748;
wire g30738;
wire g14259;
wire II37200;
wire II17662;
wire g22219;
wire g14765;
wire II40943;
wire g25181;
wire g14359;
wire II35715;
wire g26319;
wire II15949;
wire g30528;
wire g23631;
wire g21883;
wire g22552;
wire g22103;
wire g23796;
wire g23793;
wire g8978;
wire g30574;
wire g5330;
wire g16400;
wire g12215;
wire g20879;
wire g22244;
wire g30006;
wire g29498;
wire g15740;
wire g22214;
wire g28643;
wire g23261;
wire II19869;
wire g25975;
wire g28578;
wire g23674;
wire g27792;
wire g21821;
wire g28755;
wire g18329;
wire g24225;
wire g25546;
wire II27411;
wire g25952;
wire g15031;
wire g22209;
wire g10999;
wire II26980;
wire g21407;
wire II29817;
wire g24630;
wire g23203;
wire g21884;
wire g27243;
wire g24887;
wire g13982;
wire g26379;
wire g11694;
wire g18757;
wire g22001;
wire g28418;
wire II27321;
wire g26230;
wire g13375;
wire g24794;
wire g5234;
wire II39349;
wire g28087;
wire g27868;
wire II24426;
wire II39454;
wire g5924;
wire II37319;
wire g26130;
wire g13267;
wire g30806;
wire g21561;
wire II34872;
wire II30516;
wire g25081;
wire g9351;
wire II22886;
wire g22540;
wire g24465;
wire g7156;
wire g30821;
wire g23600;
wire g22140;
wire g17340;
wire g10524;
wire g16047;
wire g25640;
wire II28527;
wire g17836;
wire II25294;
wire g26892;
wire g18872;
wire g6435;
wire g11431;
wire g23607;
wire II28038;
wire II26615;
wire g27977;
wire g16287;
wire g29504;
wire g25482;
wire g16052;
wire g22746;
wire g9468;
wire g10727;
wire g20350;
wire II24346;
wire II38190;
wire II29493;
wire g22398;
wire g18277;
wire g28119;
wire g19756;
wire II32445;
wire II24656;
wire II32575;
wire g23339;
wire g29364;
wire g21133;
wire g18226;
wire g28451;
wire g22989;
wire II25540;
wire II23442;
wire g16877;
wire g29251;
wire g28703;
wire g28352;
wire g13045;
wire g28744;
wire gbuf15;
wire g10287;
wire g17092;
wire g15487;
wire II31790;
wire II30299;
wire g15759;
wire g30311;
wire g26076;
wire g12225;
wire II28137;
wire g12270;
wire II23264;
wire g26590;
wire g19573;
wire g12056;
wire II17840;
wire g17398;
wire II20386;
wire II32886;
wire g12162;
wire II29547;
wire g22759;
wire II35419;
wire II19859;
wire II32829;
wire II36432;
wire g4997;
wire II28130;
wire g15459;
wire II22983;
wire II35351;
wire g10229;
wire g20802;
wire g19262;
wire g11541;
wire g28275;
wire II15192;
wire g28153;
wire g11871;
wire g15666;
wire g19676;
wire II23619;
wire g24108;
wire g27762;
wire g26817;
wire g20700;
wire II18824;
wire g17991;
wire g19358;
wire g20594;
wire g5973;
wire II36860;
wire g26035;
wire gbuf63;
wire g13445;
wire g30001;
wire g19666;
wire g29321;
wire g6314;
wire g13059;
wire II24710;
wire g26171;
wire g22721;
wire g24429;
wire g13344;
wire II26469;
wire g27321;
wire g9092;
wire g30542;
wire II25272;
wire g17065;
wire II20339;
wire g23843;
wire g28483;
wire g20352;
wire II15942;
wire g11621;
wire g20948;
wire g8327;
wire gbuf167;
wire II28473;
wire g4067;
wire g23667;
wire g16625;
wire II24111;
wire g19672;
wire g30486;
wire g9202;
wire g26544;
wire g12318;
wire g13631;
wire g14420;
wire g28807;
wire g11102;
wire g20534;
wire g11522;
wire g10308;
wire g22470;
wire g29583;
wire g27057;
wire g15681;
wire g27986;
wire g29408;
wire g9488;
wire g23818;
wire II24603;
wire g13152;
wire g24870;
wire g27589;
wire II33488;
wire g3650;
wire gbuf5;
wire g29618;
wire g5003;
wire II32126;
wire II30979;
wire II33667;
wire g26247;
wire II16218;
wire g14747;
wire g16347;
wire II15989;
wire g10447;
wire g11910;
wire II28461;
wire g21925;
wire g19267;
wire II22563;
wire II30104;
wire g28740;
wire g24879;
wire g9776;
wire gbuf204;
wire II37590;
wire g6167;
wire g22366;
wire g25277;
wire g4095;
wire g14830;
wire g22431;
wire g15436;
wire g26137;
wire g30459;
wire g27260;
wire g27883;
wire gbuf116;
wire g29754;
wire g20775;
wire II30389;
wire g27141;
wire g10301;
wire g4240;
wire g15580;
wire g27004;
wire g27689;
wire g24544;
wire g30509;
wire II15245;
wire g23201;
wire II18369;
wire g30741;
wire g25300;
wire g11438;
wire g28606;
wire II14246;
wire II41053;
wire II33491;
wire II26931;
wire II23093;
wire g19557;
wire g14023;
wire g26574;
wire g10730;
wire g13063;
wire g12988;
wire g19888;
wire g11700;
wire g16654;
wire II40527;
wire II36718;
wire g26254;
wire g21426;
wire g5053;
wire g5854;
wire g17695;
wire g26580;
wire g5847;
wire g12097;
wire g24838;
wire II29235;
wire g17618;
wire g24860;
wire II33514;
wire g6838;
wire g9449;
wire g29084;
wire II27667;
wire g24775;
wire g12940;
wire g18949;
wire g21373;
wire g15471;
wire II38761;
wire g20506;
wire II20455;
wire g18860;
wire g13177;
wire g20347;
wire II34701;
wire g16939;
wire g23083;
wire II25071;
wire g13671;
wire g6162;
wire g15594;
wire II16703;
wire g29053;
wire g3252;
wire g8375;
wire II33723;
wire II26444;
wire g15832;
wire g13927;
wire II18362;
wire g22405;
wire g25319;
wire g11893;
wire II19657;
wire II22852;
wire g24982;
wire II36900;
wire g14796;
wire g17303;
wire g24790;
wire g4545;
wire g15335;
wire II24732;
wire g20163;
wire II31649;
wire II18133;
wire II20264;
wire g27221;
wire II35452;
wire II32480;
wire g28371;
wire g5424;
wire g29334;
wire II33655;
wire II37906;
wire g13839;
wire II18256;
wire g30396;
wire g23185;
wire g25207;
wire g4606;
wire g23585;
wire g26029;
wire g11274;
wire II35536;
wire g28642;
wire g24540;
wire g12038;
wire g29531;
wire g19108;
wire g30378;
wire g29520;
wire II21282;
wire II34857;
wire g18862;
wire g28443;
wire g10472;
wire g30581;
wire g3773;
wire g29998;
wire g14053;
wire g4332;
wire II14731;
wire II25922;
wire g19939;
wire II25740;
wire II22382;
wire II20382;
wire g19291;
wire II16209;
wire g20970;
wire II38094;
wire g29326;
wire II16476;
wire g6140;
wire g7928;
wire g15995;
wire g19901;
wire II26458;
wire II32355;
wire g19604;
wire g22282;
wire II40266;
wire g12378;
wire g16072;
wire g24332;
wire II20559;
wire g5987;
wire g22600;
wire II40589;
wire g23709;
wire II37357;
wire g6157;
wire II36132;
wire II29481;
wire II37581;
wire g23954;
wire g27827;
wire g6294;
wire II29132;
wire g10493;
wire II30407;
wire II30944;
wire g26275;
wire g3805;
wire g29355;
wire g16984;
wire g15534;
wire g24072;
wire g23219;
wire II28360;
wire g22088;
wire g17138;
wire g16998;
wire g24495;
wire II13916;
wire g11268;
wire g11963;
wire g11039;
wire g23236;
wire g11909;
wire II38074;
wire g15591;
wire II24271;
wire g23295;
wire g29091;
wire II32568;
wire g27483;
wire g21068;
wire g13167;
wire g22483;
wire g25694;
wire g20271;
wire g29244;
wire g14132;
wire II27408;
wire g4786;
wire g23561;
wire g29153;
wire g13903;
wire II33548;
wire g27565;
wire g25234;
wire II20465;
wire II33680;
wire g12699;
wire g20883;
wire II20283;
wire II20544;
wire II24319;
wire g22199;
wire g21026;
wire g16343;
wire II40949;
wire g25104;
wire g30098;
wire g27044;
wire g24043;
wire g18568;
wire g27296;
wire g25012;
wire g27338;
wire g11875;
wire g20806;
wire g8533;
wire g9584;
wire g6298;
wire g9916;
wire g14322;
wire g28654;
wire II25966;
wire g27731;
wire g30300;
wire g15219;
wire II24352;
wire g16797;
wire II38068;
wire g8676;
wire II36927;
wire g19025;
wire g12886;
wire g28342;
wire g15913;
wire g20193;
wire g7535;
wire g17802;
wire g14263;
wire g27182;
wire g28529;
wire g26803;
wire II14593;
wire g26755;
wire g12124;
wire II25940;
wire g30032;
wire g11600;
wire g30331;
wire g4967;
wire II14891;
wire II26115;
wire II41108;
wire g30226;
wire g30748;
wire g17025;
wire g19104;
wire II17059;
wire g24360;
wire g28313;
wire II16047;
wire g21590;
wire g9727;
wire g22901;
wire g20249;
wire g26047;
wire II32451;
wire g15871;
wire g10402;
wire II33297;
wire g12120;
wire g16802;
wire g11263;
wire g26490;
wire g16856;
wire g29579;
wire II31538;
wire II23824;
wire II33714;
wire II27785;
wire II32546;
wire II15230;
wire II17878;
wire g29113;
wire g9364;
wire g19316;
wire g9013;
wire g9633;
wire g26834;
wire g30493;
wire g21951;
wire g20460;
wire II34461;
wire II24703;
wire g13330;
wire g12043;
wire g30795;
wire g14381;
wire II34842;
wire II28997;
wire g4933;
wire g10570;
wire g25377;
wire g20091;
wire g27189;
wire g18023;
wire g27906;
wire gbuf144;
wire g17159;
wire g20983;
wire g26874;
wire g16218;
wire g28771;
wire g27521;
wire g25280;
wire II39460;
wire g15247;
wire g26795;
wire II40125;
wire g7754;
wire II29539;
wire g25561;
wire g23589;
wire II40176;
wire II25189;
wire g28972;
wire g30909;
wire II34392;
wire g22248;
wire g25725;
wire g28038;
wire g16722;
wire g28408;
wire II20886;
wire g29360;
wire g28843;
wire g17278;
wire g4162;
wire II20430;
wire g12235;
wire g23057;
wire g29926;
wire g25138;
wire II39002;
wire g12560;
wire II36918;
wire g7848;
wire g20472;
wire g26711;
wire g8643;
wire g10058;
wire g29396;
wire II16193;
wire g21456;
wire II13922;
wire g30505;
wire g19716;
wire II30338;
wire g24438;
wire II31928;
wire g5915;
wire II15571;
wire g17679;
wire II29333;
wire g27612;
wire g16030;
wire g9309;
wire g21448;
wire g17631;
wire g17409;
wire g21137;
wire g28054;
wire g5609;
wire g21159;
wire g23278;
wire g11686;
wire g23558;
wire II38104;
wire g19886;
wire g11462;
wire g5246;
wire g30012;
wire g28162;
wire g16181;
wire II25549;
wire II16677;
wire g21972;
wire g23243;
wire g12962;
wire g20858;
wire II27585;
wire g12339;
wire g28405;
wire II29863;
wire II21632;
wire II40901;
wire g10232;
wire g5101;
wire g20178;
wire g22693;
wire g29080;
wire II27044;
wire g5655;
wire II15277;
wire II33670;
wire g15170;
wire II27531;
wire II16163;
wire g10326;
wire II15019;
wire g8001;
wire g14139;
wire g16019;
wire g24398;
wire g27156;
wire g26651;
wire g26736;
wire g11234;
wire g7616;
wire g10709;
wire g29848;
wire II15246;
wire g25202;
wire g25411;
wire g24060;
wire gbuf126;
wire II40146;
wire II13246;
wire II15662;
wire g29096;
wire g4372;
wire g13038;
wire II27717;
wire II17300;
wire g6118;
wire g19636;
wire g24739;
wire g26718;
wire II20643;
wire g25861;
wire II35014;
wire g5774;
wire II27167;
wire g23500;
wire g29177;
wire II29271;
wire g30831;
wire II15784;
wire g23358;
wire g19723;
wire g17460;
wire II33343;
wire g16466;
wire II32309;
wire g25940;
wire II32116;
wire g23552;
wire g26570;
wire g26013;
wire II36243;
wire g18354;
wire II15932;
wire g15346;
wire g22260;
wire II14860;
wire g22299;
wire g21724;
wire g22598;
wire g23392;
wire g24557;
wire g28526;
wire g18201;
wire II27020;
wire g23691;
wire g24531;
wire II32931;
wire g19098;
wire g13422;
wire II40877;
wire II20836;
wire g16809;
wire II32719;
wire g23399;
wire g26320;
wire II18381;
wire g9806;
wire II36524;
wire g27063;
wire II13176;
wire g7745;
wire g28718;
wire g26828;
wire g24848;
wire g23538;
wire g29302;
wire g23569;
wire II25383;
wire g19280;
wire g15421;
wire g29785;
wire g11927;
wire g24239;
wire g30582;
wire II16318;
wire g22802;
wire g28291;
wire g26900;
wire II26508;
wire g25841;
wire II21838;
wire g26612;
wire g4598;
wire g11946;
wire g23210;
wire II17143;
wire g28975;
wire g25720;
wire g29619;
wire II18190;
wire II38035;
wire g12007;
wire g10045;
wire g30130;
wire II17913;
wire g17871;
wire g28363;
wire g8024;
wire g16940;
wire g21589;
wire II17637;
wire g11290;
wire g23901;
wire II18305;
wire II36663;
wire g24550;
wire II18435;
wire II39691;
wire g26262;
wire II18500;
wire g11807;
wire g29376;
wire II16328;
wire g9748;
wire g24598;
wire g18859;
wire II30626;
wire g11105;
wire g16263;
wire g11414;
wire g29857;
wire II39059;
wire g6057;
wire II36639;
wire g26634;
wire g23623;
wire g27774;
wire g23731;
wire g25266;
wire g8511;
wire g28147;
wire g10212;
wire II33249;
wire g16379;
wire g6486;
wire g28222;
wire II39255;
wire g29955;
wire g16482;
wire g11743;
wire II22536;
wire g26579;
wire g16506;
wire g4471;
wire g23134;
wire g10115;
wire g10937;
wire II33621;
wire g27172;
wire g20976;
wire g17214;
wire g25355;
wire g25461;
wire II29606;
wire g24288;
wire g12294;
wire II18470;
wire II33335;
wire II19894;
wire g8333;
wire g24872;
wire g27319;
wire g25519;
wire II27188;
wire g10834;
wire g9927;
wire II24454;
wire g28303;
wire II35527;
wire g27219;
wire g17098;
wire II15657;
wire g27710;
wire g22334;
wire g19788;
wire g8295;
wire g29835;
wire g28175;
wire g23861;
wire II37928;
wire g19228;
wire g19746;
wire g14097;
wire II33136;
wire g13228;
wire II14976;
wire II32678;
wire II32506;
wire II34479;
wire g16608;
wire g15366;
wire II27038;
wire g5813;
wire g12503;
wire g10930;
wire g27577;
wire II15856;
wire g19188;
wire g20340;
wire g19841;
wire g7957;
wire g13161;
wire g30191;
wire g5594;
wire g30714;
wire II18350;
wire g27525;
wire II16128;
wire II34363;
wire g19116;
wire g16088;
wire g24511;
wire II14675;
wire g16101;
wire II17984;
wire g26066;
wire g30984;
wire g10651;
wire II27297;
wire II40611;
wire g23283;
wire g15618;
wire g30983;
wire II31697;
wire g14374;
wire g22678;
wire g8662;
wire II34210;
wire g19203;
wire II34108;
wire g30609;
wire II30800;
wire g12830;
wire g10967;
wire g24178;
wire g30965;
wire II17892;
wire g12743;
wire II39074;
wire g17375;
wire II40560;
wire II39922;
wire g16785;
wire g20518;
wire gbuf137;
wire II21361;
wire g19651;
wire g23800;
wire g19522;
wire g14320;
wire g21803;
wire g21229;
wire g30902;
wire g26074;
wire g23212;
wire II18569;
wire g10646;
wire g19353;
wire g30665;
wire g30838;
wire g29255;
wire g8233;
wire g27673;
wire g20110;
wire g26700;
wire g21066;
wire g21034;
wire g14229;
wire g23915;
wire g21703;
wire g25539;
wire II16990;
wire g30880;
wire g3236;
wire II25240;
wire II22706;
wire g28950;
wire II28972;
wire g30264;
wire g25629;
wire g29945;
wire g26637;
wire g20481;
wire II29283;
wire g26208;
wire g13024;
wire g9320;
wire g15762;
wire II19929;
wire II18154;
wire g27437;
wire II34773;
wire II30164;
wire g10272;
wire g27613;
wire II24298;
wire g20309;
wire g19863;
wire g20387;
wire II27311;
wire g28383;
wire g5434;
wire g15307;
wire g23725;
wire g10167;
wire g25576;
wire g14329;
wire g30660;
wire g10090;
wire II14020;
wire g20446;
wire g21737;
wire g24603;
wire g22671;
wire g30552;
wire g22238;
wire g13410;
wire g26408;
wire g21104;
wire g20813;
wire g26143;
wire g30294;
wire g13415;
wire II13104;
wire g24255;
wire II33321;
wire g12853;
wire g25453;
wire g24610;
wire g5628;
wire g28795;
wire II31808;
wire g7139;
wire g27925;
wire g4501;
wire g29573;
wire g24607;
wire g27964;
wire g18820;
wire g17654;
wire II30203;
wire g10330;
wire g12890;
wire II37304;
wire g10009;
wire II40303;
wire g15046;
wire II34800;
wire g22425;
wire II36069;
wire II35092;
wire g21246;
wire g10455;
wire g16861;
wire II39393;
wire g29469;
wire II16286;
wire g9660;
wire g13077;
wire g7861;
wire g14048;
wire II37950;
wire II28218;
wire II23258;
wire g3618;
wire g18940;
wire g4584;
wire g11262;
wire g30255;
wire g11878;
wire g17795;
wire g28789;
wire g19063;
wire II40423;
wire g13516;
wire g28441;
wire II37635;
wire g19075;
wire g20637;
wire II30779;
wire g30534;
wire g4964;
wire g12191;
wire g28076;
wire g5956;
wire g17208;
wire g5199;
wire II22990;
wire g29763;
wire g6623;
wire II23133;
wire g18829;
wire II36417;
wire II15599;
wire g26699;
wire g11687;
wire II29083;
wire g27202;
wire II13140;
wire II14920;
wire II23766;
wire g13900;
wire g12651;
wire g6776;
wire II14831;
wire g16063;
wire g22079;
wire g19599;
wire g8296;
wire g7522;
wire g10605;
wire g19168;
wire g29512;
wire II36289;
wire g19662;
wire g6056;
wire g23484;
wire g18852;
wire g28018;
wire g30080;
wire gbuf218;
wire g29109;
wire g11126;
wire II26627;
wire g27209;
wire g12794;
wire g27145;
wire g10907;
wire II31195;
wire II18521;
wire g9387;
wire g10363;
wire g9669;
wire g24485;
wire g23176;
wire g25175;
wire g4757;
wire II21404;
wire II27225;
wire g29462;
wire g4418;
wire g25475;
wire II25634;
wire g18956;
wire g19976;
wire g30913;
wire g9342;
wire g13514;
wire g19837;
wire g20317;
wire g10962;
wire II35759;
wire g13125;
wire g24899;
wire II23361;
wire II18755;
wire g23118;
wire g23516;
wire II28671;
wire g10597;
wire g11518;
wire II24272;
wire g22454;
wire II28550;
wire g24579;
wire II20613;
wire II33371;
wire II16264;
wire g26129;
wire g4617;
wire II17759;
wire II25752;
wire g23852;
wire II27267;
wire g29460;
wire II30578;
wire g4797;
wire g4724;
wire g26318;
wire g19287;
wire g26829;
wire g28100;
wire g25502;
wire g12798;
wire g20722;
wire II14002;
wire g15182;
wire g23393;
wire g5824;
wire g15130;
wire g17720;
wire g20404;
wire g10588;
wire g15841;
wire g13848;
wire g19499;
wire g28941;
wire II40465;
wire g23254;
wire g11594;
wire g22836;
wire g11524;
wire II35824;
wire II33457;
wire g15825;
wire g8313;
wire g11513;
wire g5744;
wire II32726;
wire II39029;
wire II25643;
wire II39848;
wire g13585;
wire g23711;
wire g22578;
wire g19081;
wire g27561;
wire g6023;
wire II40647;
wire II38145;
wire g13192;
wire g24482;
wire g17023;
wire II30531;
wire g19764;
wire g15694;
wire g19584;
wire II25147;
wire g9264;
wire g11881;
wire g8722;
wire g13599;
wire II31109;
wire II30905;
wire II27026;
wire g20364;
wire II39359;
wire g25055;
wire g28395;
wire II33600;
wire g27546;
wire g26355;
wire gbuf78;
wire g18566;
wire II35146;
wire g18449;
wire g30463;
wire g27628;
wire II32625;
wire g29983;
wire g6635;
wire II32098;
wire g12081;
wire g30121;
wire g20414;
wire g28691;
wire g16106;
wire II30332;
wire II30911;
wire g23159;
wire g22271;
wire II37008;
wire g14194;
wire g28948;
wire g22618;
wire g17540;
wire g30020;
wire g10104;
wire g28269;
wire g30864;
wire g23221;
wire g10173;
wire II26926;
wire II22163;
wire g17775;
wire II24306;
wire g24822;
wire g3957;
wire II24476;
wire g15093;
wire g18543;
wire g25060;
wire II31793;
wire g25669;
wire g29612;
wire g29483;
wire II21881;
wire g13031;
wire II21761;
wire g12871;
wire II13421;
wire g10375;
wire g22149;
wire g23340;
wire g18844;
wire g19167;
wire g15605;
wire g16311;
wire g11945;
wire g20841;
wire II13478;
wire II15445;
wire g30350;
wire g15145;
wire g21385;
wire g13855;
wire g24524;
wire II27218;
wire g5950;
wire II28103;
wire g9726;
wire II17649;
wire g24283;
wire g27701;
wire g20897;
wire g10369;
wire g13676;
wire g30940;
wire II26317;
wire g16141;
wire II37122;
wire g18602;
wire g4760;
wire II24186;
wire g12299;
wire g19830;
wire g18637;
wire II23932;
wire g29913;
wire g10887;
wire g16425;
wire g26344;
wire g10480;
wire g23163;
wire g24570;
wire g20337;
wire II30380;
wire II22775;
wire II34132;
wire g30519;
wire g30500;
wire g19252;
wire II37143;
wire g30063;
wire g27506;
wire II26123;
wire g14106;
wire g21844;
wire g27909;
wire II20132;
wire g20150;
wire g18509;
wire g13818;
wire g11246;
wire II30311;
wire II30353;
wire II24596;
wire g12547;
wire II28506;
wire g8303;
wire g9888;
wire II36060;
wire g21188;
wire II26999;
wire II39825;
wire II29641;
wire g27579;
wire g20684;
wire g21825;
wire g8898;
wire g5768;
wire II28781;
wire g12783;
wire g24247;
wire g28172;
wire II39806;
wire II25573;
wire II39832;
wire g5684;
wire g27000;
wire g25069;
wire II16835;
wire g15725;
wire II35768;
wire g15797;
wire g14041;
wire g5067;
wire g20466;
wire g24503;
wire g13434;
wire g14514;
wire II32616;
wire g24420;
wire g4310;
wire g15962;
wire g20250;
wire II38440;
wire g26748;
wire II40188;
wire g18934;
wire g28461;
wire g5785;
wire g19942;
wire g12444;
wire g13132;
wire g16905;
wire g27583;
wire II28557;
wire II28966;
wire g27022;
wire g6215;
wire g23156;
wire g10296;
wire g25242;
wire II30329;
wire g29227;
wire II32499;
wire g12273;
wire II38698;
wire II40817;
wire II35904;
wire g22547;
wire g11202;
wire g29655;
wire II31835;
wire g21577;
wire II35506;
wire g13274;
wire g30742;
wire g24241;
wire g27395;
wire g22581;
wire II22503;
wire II34421;
wire g5293;
wire g30722;
wire g21685;
wire g22806;
wire g13644;
wire g26859;
wire II18593;
wire g5806;
wire II24166;
wire g9107;
wire II24053;
wire g25557;
wire II14384;
wire II13971;
wire g30394;
wire g22038;
wire II37312;
wire g23003;
wire g16656;
wire g23950;
wire II33954;
wire g8798;
wire g28116;
wire g23894;
wire g13458;
wire g29183;
wire II13601;
wire II27949;
wire g18688;
wire g26661;
wire g23572;
wire g26250;
wire II38184;
wire g20994;
wire g21207;
wire g20087;
wire II21476;
wire g11709;
wire g29471;
wire g13040;
wire II23374;
wire g28158;
wire II24408;
wire g10262;
wire II25054;
wire g16830;
wire II27388;
wire g5704;
wire g27911;
wire g22917;
wire g10468;
wire g7632;
wire g16057;
wire g25162;
wire g21428;
wire II29177;
wire g21721;
wire g20991;
wire g11182;
wire g23021;
wire g9114;
wire g17649;
wire II30881;
wire g27446;
wire g8778;
wire g19825;
wire g25225;
wire g22382;
wire g13493;
wire II36114;
wire g25895;
wire g24583;
wire g27165;
wire g8524;
wire g21508;
wire g21182;
wire g8820;
wire II33999;
wire g8529;
wire II34866;
wire II23395;
wire g25985;
wire g27655;
wire g19615;
wire II34059;
wire g25931;
wire g24567;
wire g26325;
wire g22643;
wire g29701;
wire II26006;
wire g17719;
wire II18378;
wire g27970;
wire II18423;
wire g4453;
wire g13249;
wire g21695;
wire II13745;
wire II21644;
wire g10413;
wire g11783;
wire g17246;
wire II21435;
wire II32181;
wire g28288;
wire II22318;
wire gbuf191;
wire gbuf166;
wire g17193;
wire II15645;
wire II30239;
wire II26407;
wire g12600;
wire II16159;
wire g27062;
wire g21872;
wire g23497;
wire g13837;
wire g15839;
wire II38272;
wire II36687;
wire g12981;
wire II31811;
wire g10145;
wire g19697;
wire g14423;
wire g10038;
wire g30499;
wire g15391;
wire g29261;
wire II38653;
wire g23080;
wire g16535;
wire g20578;
wire g4489;
wire g28056;
wire g27029;
wire g27971;
wire g5618;
wire g13703;
wire II28335;
wire g21263;
wire g15625;
wire g20427;
wire II20376;
wire II28432;
wire g19272;
wire g9288;
wire g4326;
wire II24466;
wire g29409;
wire g12820;
wire g12435;
wire g29222;
wire g12204;
wire II22136;
wire g22975;
wire g16820;
wire II21583;
wire g27672;
wire g10473;
wire g10394;
wire g12022;
wire g14092;
wire g18059;
wire g24122;
wire g26559;
wire II31077;
wire II32411;
wire g29190;
wire g24611;
wire g5200;
wire II32559;
wire g18084;
wire g24784;
wire g21085;
wire g16686;
wire g21352;
wire g30675;
wire g23097;
wire g15650;
wire II25018;
wire g23324;
wire g13407;
wire g21141;
wire II25690;
wire g25255;
wire g29127;
wire g30852;
wire g6513;
wire II28515;
wire II33157;
wire II40498;
wire II30679;
wire g19733;
wire g16451;
wire g29371;
wire II24459;
wire II26996;
wire g16444;
wire g17063;
wire g19414;
wire g17979;
wire g9871;
wire g11644;
wire g12938;
wire g12107;
wire II32709;
wire g5909;
wire g13612;
wire g26081;
wire g16220;
wire g8860;
wire g23223;
wire g24889;
wire II19160;
wire g23172;
wire g21346;
wire g5641;
wire II36963;
wire II37602;
wire g10481;
wire g10469;
wire II38817;
wire g13475;
wire g15415;
wire g20669;
wire g20022;
wire II38136;
wire g13609;
wire g4567;
wire g9670;
wire II24247;
wire g30233;
wire g13396;
wire g15750;
wire II25617;
wire g27356;
wire g19430;
wire g28820;
wire II16972;
wire g13054;
wire g22683;
wire II31817;
wire g5837;
wire g29438;
wire g19182;
wire g26925;
wire g12267;
wire II25377;
wire g26741;
wire II30470;
wire g23103;
wire g8605;
wire g20160;
wire g22707;
wire II32057;
wire g27989;
wire g10987;
wire g27277;
wire g9073;
wire g19040;
wire g23141;
wire II36330;
wire g22090;
wire g11530;
wire II24634;
wire g9212;
wire II18405;
wire g16241;
wire II28190;
wire g5078;
wire g23665;
wire g11425;
wire g25708;
wire II27689;
wire g22922;
wire g23040;
wire g29632;
wire g18717;
wire II16234;
wire g29778;
wire II31112;
wire g12174;
wire g18370;
wire g25938;
wire II24125;
wire g24296;
wire g27084;
wire g10206;
wire g24321;
wire g20934;
wire g20564;
wire II23466;
wire g25153;
wire g4295;
wire II39148;
wire g26589;
wire g11769;
wire g4204;
wire g19208;
wire g26163;
wire g22666;
wire II26777;
wire g24265;
wire g17527;
wire gbuf94;
wire g30759;
wire g13914;
wire II33573;
wire g4737;
wire g20343;
wire II21677;
wire g21758;
wire II33624;
wire g11918;
wire g27741;
wire g21688;
wire g21762;
wire gbuf133;
wire g30972;
wire g15311;
wire g25553;
wire g22656;
wire g20115;
wire g17685;
wire g26470;
wire g27248;
wire g24799;
wire g21328;
wire g9647;
wire g28499;
wire g10533;
wire g26001;
wire g8397;
wire g22162;
wire g21879;
wire g29199;
wire g16002;
wire g16596;
wire II23553;
wire g17445;
wire g25773;
wire g15802;
wire g15761;
wire g20585;
wire II40044;
wire II34099;
wire II34806;
wire II15967;
wire II16776;
wire g17517;
wire g25490;
wire g28474;
wire II34821;
wire g10380;
wire g24092;
wire g5071;
wire g26405;
wire g11002;
wire g10591;
wire II14668;
wire gbuf148;
wire II28447;
wire g20106;
wire II37968;
wire II22028;
wire g9534;
wire g5928;
wire g14079;
wire g7751;
wire g24270;
wire g22235;
wire II38491;
wire II29462;
wire g22714;
wire g29644;
wire g7772;
wire II18725;
wire II13501;
wire g29793;
wire g17171;
wire gbuf86;
wire g25020;
wire g15951;
wire g24229;
wire II16881;
wire g26479;
wire II37062;
wire g30661;
wire g29809;
wire g20216;
wire g5033;
wire g19324;
wire g3999;
wire g27175;
wire II35994;
wire g16120;
wire g10108;
wire g21689;
wire g19417;
wire g25995;
wire g16566;
wire II14416;
wire II36264;
wire II36527;
wire II38656;
wire II16024;
wire g23939;
wire g8612;
wire g22526;
wire g23638;
wire II41044;
wire g24923;
wire II39154;
wire g12519;
wire II14934;
wire g22205;
wire II18857;
wire II31165;
wire g6707;
wire g15021;
wire g13480;
wire g30399;
wire g28457;
wire g27861;
wire g16321;
wire II40673;
wire g19467;
wire g26039;
wire g11176;
wire g28450;
wire g4656;
wire g11291;
wire g5708;
wire g27078;
wire II24214;
wire g12434;
wire II21730;
wire g18547;
wire g14360;
wire g7465;
wire g22098;
wire g25221;
wire II18473;
wire g21075;
wire g7875;
wire II28351;
wire II38229;
wire g8655;
wire g27233;
wire II18707;
wire g7823;
wire II34172;
wire II34839;
wire g6153;
wire g16629;
wire g10890;
wire II24071;
wire g20623;
wire II32596;
wire II37569;
wire g20289;
wire g15828;
wire g8774;
wire g30825;
wire g9747;
wire g10066;
wire II36450;
wire g7792;
wire g26560;
wire g20378;
wire II40197;
wire g26024;
wire g29073;
wire g15283;
wire g27159;
wire II38391;
wire g13623;
wire II38804;
wire II34671;
wire II19602;
wire II19455;
wire g26668;
wire II38032;
wire g21283;
wire g27688;
wire II35123;
wire g29163;
wire gbuf214;
wire g23821;
wire g7259;
wire II36302;
wire g26549;
wire II39331;
wire II18344;
wire II25731;
wire g16994;
wire gbuf47;
wire g10549;
wire g22864;
wire II37917;
wire II31826;
wire g19455;
wire g27790;
wire g27194;
wire g24853;
wire g15615;
wire g12181;
wire g21323;
wire g13206;
wire g16433;
wire II24415;
wire g27387;
wire g5860;
wire g21360;
wire g29278;
wire g24788;
wire g30895;
wire g25458;
wire g13223;
wire g20398;
wire g28837;
wire g26485;
wire g25077;
wire g12250;
wire g11148;
wire II35953;
wire g16262;
wire g17573;
wire II22545;
wire g7303;
wire g13146;
wire II24565;
wire g11539;
wire g9025;
wire g17655;
wire g22081;
wire g8626;
wire g13116;
wire g23120;
wire g25103;
wire II23673;
wire g15356;
wire g15670;
wire g13361;
wire g22173;
wire g30950;
wire II33816;
wire g6038;
wire g29959;
wire g6288;
wire g13255;
wire g19770;
wire II36666;
wire II18259;
wire g30989;
wire II19631;
wire II32588;
wire g13487;
wire g11637;
wire g22791;
wire II15671;
wire g30365;
wire g21019;
wire g28715;
wire g10566;
wire g19101;
wire II36102;
wire g4217;
wire g26175;
wire II18107;
wire g14207;
wire II21488;
wire II24236;
wire g18825;
wire II27005;
wire g5886;
wire II32970;
wire g5639;
wire g26794;
wire g29667;
wire g29235;
wire g27470;
wire g20187;
wire g25050;
wire II18097;
wire g3940;
wire g5793;
wire g27875;
wire g8236;
wire g30309;
wire g29205;
wire g22046;
wire g5550;
wire g12239;
wire II35053;
wire g29292;
wire g10613;
wire g3942;
wire g17927;
wire g23873;
wire g15290;
wire II16006;
wire g29658;
wire II40829;
wire g26971;
wire g29026;
wire g28490;
wire II30965;
wire g11364;
wire II27382;
wire g20703;
wire II38841;
wire g24355;
wire g20441;
wire g26096;
wire g11209;
wire g6443;
wire g23127;
wire g25418;
wire II18662;
wire g27991;
wire g23525;
wire g19263;
wire g4133;
wire g21901;
wire g23539;
wire g11309;
wire II20547;
wire g30953;
wire II40143;
wire g15661;
wire g30034;
wire II30728;
wire g8147;
wire g27518;
wire g11891;
wire II29336;
wire g13572;
wire g25755;
wire g28832;
wire II33408;
wire g27308;
wire II18746;
wire g24436;
wire g30554;
wire g28955;
wire g25044;
wire g8439;
wire II36721;
wire g26333;
wire g14153;
wire g30472;
wire II13968;
wire g28479;
wire g5132;
wire II25882;
wire g24728;
wire g23899;
wire g11984;
wire II39014;
wire g29802;
wire g10121;
wire g16814;
wire II34143;
wire g26385;
wire g21963;
wire II24502;
wire II25153;
wire g11475;
wire g26269;
wire g24975;
wire g23629;
wire II31715;
wire II41141;
wire g8089;
wire g10943;
wire g19300;
wire g19817;
wire g20936;
wire g20962;
wire g29218;
wire g21128;
wire gbuf97;
wire g21856;
wire g26059;
wire g15235;
wire g24309;
wire g19034;
wire II40075;
wire II27065;
wire g26294;
wire g24752;
wire g21311;
wire g15464;
wire g26812;
wire II14766;
wire g7574;
wire II29383;
wire II27537;
wire g23409;
wire g22733;
wire g23402;
wire g20290;
wire g30389;
wire g26978;
wire II40712;
wire g30093;
wire g18611;
wire g30221;
wire g18806;
wire g17635;
wire g21482;
wire II28374;
wire g30324;
wire g23148;
wire g8466;
wire II23941;
wire g18108;
wire II38471;
wire II33640;
wire g24344;
wire II25168;
wire g19589;
wire g10432;
wire g17272;
wire II30786;
wire II40967;
wire g9140;
wire g19872;
wire g16020;
wire g10876;
wire II28271;
wire II15183;
wire II38107;
wire II14091;
wire g26493;
wire g28676;
wire g26867;
wire g29975;
wire g18014;
wire g18405;
wire II29180;
wire g23460;
wire g26725;
wire g20493;
wire g19925;
wire g16650;
wire g9131;
wire g20306;
wire II34241;
wire II27056;
wire g27569;
wire II22283;
wire g30490;
wire g15374;
wire g23622;
wire g18707;
wire II40658;
wire g27135;
wire g18363;
wire g28583;
wire g30402;
wire II37641;
wire g11563;
wire g23316;
wire II19642;
wire g20830;
wire g13308;
wire g24769;
wire g18789;
wire II31748;
wire g8812;
wire g21092;
wire II29715;
wire g13028;
wire II16694;
wire g5613;
wire g21050;
wire g8649;
wire g22787;
wire g20925;
wire g28712;
wire II39785;
wire II39585;
wire g10974;
wire g26967;
wire g28554;
wire g25176;
wire g26994;
wire g3246;
wire g15260;
wire II17743;
wire g12705;
wire g27681;
wire II36393;
wire II31541;
wire g30506;
wire II16196;
wire g24500;
wire g28629;
wire II29906;
wire g8979;
wire g30412;
wire g7619;
wire g30466;
wire II37002;
wire g27344;
wire g19321;
wire g23126;
wire g11788;
wire g10735;
wire g18296;
wire g16848;
wire g11532;
wire g30819;
wire g21345;
wire g30107;
wire g4272;
wire g12040;
wire g23464;
wire g29179;
wire g18900;
wire II31943;
wire g30380;
wire II26365;
wire II33472;
wire II14709;
wire II30931;
wire g30343;
wire g29315;
wire g10439;
wire g19576;
wire g29925;
wire g25609;
wire g26229;
wire II15190;
wire g4041;
wire g22066;
wire g20299;
wire g30958;
wire g12941;
wire g10399;
wire g16614;
wire II38662;
wire g22843;
wire g11957;
wire g21715;
wire II26645;
wire g26673;
wire II35945;
wire g27690;
wire g8878;
wire g29537;
wire II36969;
wire g28759;
wire II29536;
wire g4827;
wire II19797;
wire g15831;
wire II36659;
wire II28991;
wire g8868;
wire g21748;
wire g1248;
wire g16006;
wire g29038;
wire II27285;
wire II15535;
wire g25351;
wire g23119;
wire II19030;
wire g22725;
wire g16492;
wire g21413;
wire II38379;
wire g28469;
wire g24949;
wire g8505;
wire g16825;
wire II27779;
wire g26569;
wire g29141;
wire II31445;
wire II37956;
wire g24641;
wire g21948;
wire g25287;
wire g30510;
wire g16384;
wire g20631;
wire g17937;
wire g17761;
wire II17981;
wire II13504;
wire g28024;
wire g11527;
wire II16357;
wire II34860;
wire g12647;
wire II30504;
wire g29196;
wire g7573;
wire g18782;
wire g30761;
wire II19618;
wire g13974;
wire g10478;
wire II23636;
wire II18302;
wire g22181;
wire g12155;
wire g7532;
wire II15454;
wire II25253;
wire g16967;
wire g9661;
wire g22188;
wire g22223;
wire g12880;
wire g23714;
wire g28216;
wire g15032;
wire g23543;
wire g20566;
wire g8908;
wire g26234;
wire g9481;
wire II21615;
wire g10745;
wire g4465;
wire g17429;
wire g22596;
wire g5664;
wire g5960;
wire g20826;
wire g26652;
wire II39919;
wire g11973;
wire II33385;
wire II20640;
wire g26018;
wire g24400;
wire g11138;
wire g27431;
wire II16438;
wire g21053;
wire g25027;
wire g30390;
wire II16107;
wire II13892;
wire g28853;
wire g26365;
wire g11934;
wire g13548;
wire g19919;
wire II34971;
wire g9734;
wire g14238;
wire g10670;
wire g18074;
wire g23532;
wire g17209;
wire II35485;
wire g12538;
wire g23683;
wire II40709;
wire II27300;
wire II38396;
wire II26085;
wire g13189;
wire g17202;
wire g23145;
wire g21597;
wire g8388;
wire g25121;
wire gbuf101;
wire g13530;
wire II31152;
wire g23448;
wire g30768;
wire II33649;
wire g25237;
wire g8839;
wire g16395;
wire g21435;
wire g29561;
wire II15546;
wire g9057;
wire g19621;
wire g25618;
wire g29934;
wire g11958;
wire II40691;
wire II37280;
wire II37074;
wire II38722;
wire g10452;
wire g29986;
wire II16335;
wire g11949;
wire II36493;
wire g8714;
wire g16847;
wire g27097;
wire g11435;
wire g26567;
wire g4015;
wire g29456;
wire g24293;
wire g15220;
wire g21340;
wire g25826;
wire g30871;
wire g21953;
wire g18325;
wire g28082;
wire g11404;
wire g10063;
wire g20422;
wire g17167;
wire g23728;
wire g12075;
wire g21173;
wire g5064;
wire II28123;
wire II33662;
wire g26340;
wire g28166;
wire g4905;
wire g29280;
wire II38851;
wire g13529;
wire II23029;
wire g15755;
wire II18375;
wire g5859;
wire g10520;
wire gbuf99;
wire g28244;
wire g8573;
wire g19354;
wire g21316;
wire g26941;
wire II24263;
wire II38857;
wire g23922;
wire g17716;
wire g22607;
wire II13101;
wire g21887;
wire g27089;
wire g24263;
wire g11999;
wire g26025;
wire g27312;
wire g23604;
wire g4101;
wire g23309;
wire g20940;
wire g4541;
wire g26681;
wire g21377;
wire g19309;
wire g22985;
wire II14778;
wire g6912;
wire g26896;
wire g21293;
wire g17366;
wire g19931;
wire II24124;
wire g28782;
wire g11579;
wire g28334;
wire g15898;
wire g24779;
wire II14249;
wire II37134;
wire II19307;
wire g15807;
wire g4003;
wire g19812;
wire g18221;
wire II30803;
wire g29325;
wire g16895;
wire II25283;
wire g26763;
wire II28464;
wire g13285;
wire g22669;
wire g22004;
wire g26188;
wire II27116;
wire g18618;
wire g28748;
wire g4928;
wire g10305;
wire g30089;
wire g30565;
wire g5238;
wire g13049;
wire g10227;
wire g25505;
wire g7153;
wire g11627;
wire g11896;
wire II36996;
wire g11582;
wire II36272;
wire g19546;
wire g24590;
wire g24676;
wire g8252;
wire g29404;
wire II41050;
wire g10867;
wire g18667;
wire II24608;
wire g20138;
wire g12454;
wire g30315;
wire II28741;
wire g26556;
wire g18063;
wire g23847;
wire g11967;
wire II30236;
wire g4632;
wire g5751;
wire g17551;
wire II24916;
wire g22144;
wire II37032;
wire g25144;
wire g19046;
wire g25257;
wire g17947;
wire g8761;
wire g15756;
wire g5903;
wire II18620;
wire g20356;
wire II29936;
wire g22742;
wire II38875;
wire gbuf67;
wire g10574;
wire g3677;
wire II15304;
wire g8911;
wire g20805;
wire g24460;
wire II30594;
wire II30401;
wire g19161;
wire g27365;
wire II31619;
wire gbuf196;
wire g29759;
wire g25065;
wire gbuf11;
wire g16133;
wire g24104;
wire g4486;
wire g9521;
wire g18753;
wire g27215;
wire g9463;
wire g14464;
wire g21817;
wire II37179;
wire g18491;
wire g6166;
wire II33888;
wire g19771;
wire g7265;
wire g30966;
wire g27005;
wire II35079;
wire g17912;
wire g11778;
wire II24389;
wire g22342;
wire g29689;
wire g10996;
wire II30894;
wire g11770;
wire g17384;
wire g21541;
wire g24864;
wire g4203;
wire g12148;
wire II29927;
wire g29063;
wire g29382;
wire g5118;
wire g23046;
wire II23115;
wire g20622;
wire g12415;
wire g22935;
wire g25304;
wire g26414;
wire II33517;
wire g24425;
wire g27017;
wire g25430;
wire g4185;
wire g29994;
wire g24638;
wire g25678;
wire g27053;
wire g26259;
wire g6783;
wire II17670;
wire g25204;
wire II31832;
wire g29905;
wire g22061;
wire g26895;
wire II18524;
wire g27397;
wire g19660;
wire II38701;
wire g20985;
wire g16211;
wire g26979;
wire gbuf31;
wire g19914;
wire II24950;
wire g16644;
wire g22362;
wire II37494;
wire II23806;
wire g23153;
wire II18787;
wire II16747;
wire g27742;
wire II23457;
wire g23181;
wire g11281;
wire g18107;
wire g25915;
wire g11837;
wire g20050;
wire g28636;
wire g28279;
wire II31454;
wire g11703;
wire II33495;
wire II31763;
wire II36808;
wire g30850;
wire g21162;
wire g11598;
wire g28487;
wire g23592;
wire g11459;
wire g23094;
wire g27289;
wire II17910;
wire g24875;
wire g10261;
wire II32320;
wire g6448;
wire g27355;
wire g18526;
wire g19564;
wire II22952;
wire g29548;
wire g29966;
wire g7459;
wire g9083;
wire g21422;
wire g24415;
wire g5851;
wire II35021;
wire g18977;
wire II17816;
wire g29329;
wire II32346;
wire g29840;
wire g13878;
wire II31127;
wire g25980;
wire g29119;
wire g5716;
wire g13873;
wire II29613;
wire g17116;
wire g5705;
wire g11914;
wire g19500;
wire II18943;
wire g20502;
wire II29360;
wire g5651;
wire gbuf112;
wire g23300;
wire g28669;
wire II39930;
wire g13055;
wire g27048;
wire g15019;
wire II18204;
wire g9891;
wire II24743;
wire g30869;
wire g17507;
wire g29529;
wire II18777;
wire g30844;
wire g29535;
wire II16876;
wire g19347;
wire II18566;
wire g10014;
wire g9922;
wire g13934;
wire g4945;
wire II33659;
wire g17393;
wire II38408;
wire g28894;
wire g12034;
wire g29607;
wire g25315;
wire g3235;
wire g6430;
wire g3243;
wire g23505;
wire g29410;
wire II13128;
wire g13464;
wire g13632;
wire g23315;
wire II36123;
wire g20738;
wire g9591;
wire g11591;
wire g19688;
wire g26531;
wire g7607;
wire g20679;
wire g12863;
wire g20457;
wire II19628;
wire g24055;
wire g24644;
wire g13600;
wire II31655;
wire II19105;
wire g28962;
wire g13881;
wire II30525;
wire g29264;
wire g26070;
wire g11589;
wire g16770;
wire g30919;
wire II33434;
wire g8406;
wire II16156;
wire g4415;
wire II30763;
wire g21789;
wire g18874;
wire g22231;
wire gbuf189;
wire g10289;
wire g24507;
wire g15744;
wire II17060;
wire g15784;
wire g18952;
wire II27095;
wire g22182;
wire g30539;
wire g20145;
wire g25184;
wire g12996;
wire g25179;
wire g30929;
wire II24061;
wire g27717;
wire II31290;
wire g20012;
wire II16120;
wire g18832;
wire g28265;
wire g9794;
wire g26113;
wire g19213;
wire g30071;
wire g6641;
wire g9762;
wire II39913;
wire g23972;
wire g7898;
wire g22307;
wire g23677;
wire g25372;
wire g20554;
wire g20016;
wire g17080;
wire g21996;
wire g29726;
wire II18329;
wire g18867;
wire g22628;
wire g10556;
wire g21195;
wire g15845;
wire g30935;
wire g5213;
wire g19705;
wire g24835;
wire g8958;
wire g20297;
wire II37273;
wire g24212;
wire II34114;
wire g21397;
wire g30687;
wire g13958;
wire g16170;
wire g26196;
wire g21009;
wire g9905;
wire II26340;
wire g8843;
wire II23742;
wire g26539;
wire g5879;
wire g14107;
wire g8723;
wire g25361;
wire II29951;
wire g13120;
wire g21628;
wire II17070;
wire g11712;
wire g19767;
wire g30455;
wire g12913;
wire g23024;
wire g18246;
wire g18805;
wire g18985;
wire g18586;
wire g27113;
wire g8414;
wire g16356;
wire g11225;
wire g29131;
wire g22613;
wire II37863;
wire g5921;
wire II18810;
wire g20324;
wire g30461;
wire g25954;
wire g23797;
wire g30653;
wire g25437;
wire II36621;
wire gbuf151;
wire g8763;
wire g11826;
wire g19780;
wire g30064;
wire II35731;
wire g7337;
wire g13791;
wire g6204;
wire g22992;
wire g24457;
wire g27096;
wire g10372;
wire g16236;
wire II37170;
wire II28988;
wire II23173;
wire g13455;
wire g6894;
wire II29465;
wire g24454;
wire g22125;
wire g26758;
wire II21888;
wire g25347;
wire II16344;
wire II29116;
wire II15478;
wire g16693;
wire II24077;
wire g14960;
wire g28121;
wire II20328;
wire II27355;
wire g30680;
wire g23031;
wire II14066;
wire g18921;
wire II28143;
wire g30878;
wire g5999;
wire g8544;
wire g19259;
wire g19712;
wire g9752;
wire g6177;
wire g29546;
wire g22633;
wire II23242;
wire g13168;
wire g13441;
wire II17483;
wire II15696;
wire g19244;
wire II18043;
wire II34668;
wire g9146;
wire II18295;
wire g11853;
wire g19693;
wire II40979;
wire g6131;
wire g17155;
wire g10787;
wire g30694;
wire g26841;
wire II40627;
wire II30660;
wire g7527;
wire g13582;
wire II27032;
wire g18237;
wire II23020;
wire g16456;
wire II21321;
wire g20913;
wire g23483;
wire g18826;
wire g25294;
wire II25562;
wire g12209;
wire II40694;
wire g5870;
wire g30546;
wire g16640;
wire g19011;
wire g22737;
wire g26140;
wire g24627;
wire g5342;
wire II29945;
wire II24758;
wire II13134;
wire g25340;
wire g12325;
wire g15454;
wire g30922;
wire g27935;
wire g13824;
wire g15540;
wire g5473;
wire g6193;
wire g30143;
wire g12061;
wire g6062;
wire g25009;
wire g24163;
wire g4347;
wire g18147;
wire g14355;
wire II23658;
wire g17056;
wire g27549;
wire g19386;
wire II40584;
wire II36521;
wire II27215;
wire II21374;
wire g20891;
wire II19271;
wire II23392;
wire g22777;
wire g22762;
wire II31787;
wire g24313;
wire g8974;
wire g26105;
wire g30586;
wire II21949;
wire II38241;
wire g22112;
wire g18090;
wire g24209;
wire g15096;
wire g5257;
wire g27390;
wire II34189;
wire g17604;
wire g25385;
wire g5867;
wire g22847;
wire g20604;
wire g10889;
wire g21895;
wire II16562;
wire g13501;
wire II35428;
wire II15879;
wire II20622;
wire g29447;
wire g24284;
wire g30118;
wire II20365;
wire g21370;
wire g24818;
wire g4692;
wire g29454;
wire g20373;
wire g18835;
wire II27695;
wire g29677;
wire g20403;
wire g17224;
wire g30048;
wire g7622;
wire g11940;
wire g27226;
wire g10801;
wire g9139;
wire II35863;
wire g11519;
wire g6908;
wire II16138;
wire g14316;
wire g27769;
wire II15909;
wire g16301;
wire g25869;
wire g8160;
wire g9063;
wire II24300;
wire II31901;
wire II29687;
wire II23929;
wire g30524;
wire g7993;
wire g7976;
wire g15537;
wire g22295;
wire g22016;
wire g13318;
wire g29297;
wire g19920;
wire g23069;
wire g9932;
wire g30734;
wire g24813;
wire II13575;
wire g20039;
wire g19853;
wire II17869;
wire g16404;
wire g26617;
wire II33330;
wire g24844;
wire II24507;
wire g19453;
wire g22753;
wire g25945;
wire g30971;
wire g23138;
wire II29550;
wire g28057;
wire g10276;
wire g28610;
wire g17259;
wire g21593;
wire II30383;
wire g19728;
wire II38650;
wire g13245;
wire g28050;
wire g19791;
wire II24235;
wire g19009;
wire II40230;
wire g20955;
wire g19286;
wire g10103;
wire g10446;
wire g29606;
wire II32487;
wire g25263;
wire g25167;
wire g21179;
wire II40113;
wire II28482;
wire g30884;
wire g9341;
wire II34395;
wire g16486;
wire g12744;
wire g28115;
wire g12232;
wire g5626;
wire g24142;
wire g16253;
wire g3462;
wire g29161;
wire g23152;
wire II20556;
wire g8499;
wire g30060;
wire g15409;
wire g16884;
wire II40051;
wire g26217;
wire II35095;
wire g5243;
wire II35341;
wire g20760;
wire g23434;
wire g30134;
wire II39035;
wire g13425;
wire g13451;
wire g30711;
wire g10797;
wire g29306;
wire g23287;
wire g17236;
wire II37400;
wire g5385;
wire g6897;
wire g5438;
wire g9323;
wire g29399;
wire II16779;
wire II30059;
wire g10094;
wire g19284;
wire g4474;
wire II24662;
wire g23168;
wire g23471;
wire g21415;
wire g26551;
wire g27529;
wire g16367;
wire g26290;
wire g13124;
wire g13834;
wire II34776;
wire g20407;
wire g20581;
wire g22825;
wire g5507;
wire g20652;
wire II25899;
wire g11774;
wire g15679;
wire g11921;
wire g19578;
wire g28070;
wire g23828;
wire g8209;
wire g15177;
wire II36507;
wire g27231;
wire g17228;
wire II39083;
wire II18411;
wire g23311;
wire g8700;
wire g27754;
wire II20305;
wire II25702;
wire g19550;
wire II33260;
wire g25247;
wire II19937;
wire II35043;
wire g21791;
wire g20969;
wire g29990;
wire II35364;
wire g6216;
wire g24749;
wire II39020;
wire II13950;
wire g24554;
wire g15545;
wire II31736;
wire g13142;
wire g11063;
wire g12362;
wire II30476;
wire g15426;
wire g12858;
wire g30798;
wire g5114;
wire g27892;
wire g19656;
wire g23943;
wire g21573;
wire g11552;
wire g23415;
wire g24476;
wire g5816;
wire II21691;
wire g23786;
wire g29372;
wire g9102;
wire g24079;
wire g27050;
wire g28226;
wire g22729;
wire g19224;
wire g15161;
wire g13546;
wire g8971;
wire g25218;
wire g22274;
wire II23009;
wire g4424;
wire g29946;
wire g30195;
wire g23735;
wire II40317;
wire g28751;
wire II32677;
wire g4441;
wire g9497;
wire II17798;
wire g25514;
wire II18280;
wire g4868;
wire II33396;
wire g16013;
wire gbuf209;
wire g27573;
wire g11798;
wire II34794;
wire II41138;
wire g5899;
wire g15765;
wire g20665;
wire g7953;
wire II28027;
wire g29979;
wire g28331;
wire g24515;
wire II16507;
wire II29591;
wire II38214;
wire gbuf62;
wire g19779;
wire g22484;
wire g5362;
wire g10459;
wire g11421;
wire II29700;
wire g15942;
wire g24499;
wire g22837;
wire g16111;
wire II22444;
wire g20485;
wire g26850;
wire g20902;
wire g15821;
wire II28789;
wire g8492;
wire g20081;
wire g15043;
wire II16611;
wire g18670;
wire g22722;
wire g10542;
wire g28148;
wire g17378;
wire g22566;
wire g23376;
wire II14993;
wire II18281;
wire g24381;
wire g25723;
wire II15610;
wire g28296;
wire g29559;
wire g20783;
wire g21809;
wire II30648;
wire g23565;
wire g20501;
wire g25797;
wire g24001;
wire g25272;
wire II29445;
wire g23748;
wire g4444;
wire g18814;
wire II25664;
wire g25155;
wire g21225;
wire g28307;
wire g3900;
wire g12522;
wire g10640;
wire g21867;
wire II36761;
wire g28043;
wire g21027;
wire II25001;
wire g3997;
wire g28096;
wire g29698;
wire g18910;
wire II23225;
wire g22055;
wire g8568;
wire g18654;
wire g21337;
wire g21899;
wire II32461;
wire g21307;
wire II34068;
wire g25403;
wire II19753;
wire II19374;
wire g17020;
wire g30291;
wire g27543;
wire g30298;
wire g9067;
wire g16559;
wire II22789;
wire g4269;
wire g17288;
wire g12431;
wire II32898;
wire II35799;
wire II32835;
wire g15493;
wire g11804;
wire g22996;
wire g15766;
wire II16931;
wire g23419;
wire II38898;
wire g28799;
wire g30777;
wire g16448;
wire g19144;
wire g29659;
wire g14233;
wire g24928;
wire g17217;
wire g29950;
wire II30365;
wire g30980;
wire g22768;
wire g22799;
wire g26704;
wire g5597;
wire g29821;
wire II32267;
wire g17799;
wire II35524;
wire g30745;
wire g17807;
wire II26690;
wire II40206;
wire II18287;
wire g19164;
wire g21911;
wire g27811;
wire g27968;
wire g15440;
wire II24361;
wire II16552;
wire g13395;
wire g23016;
wire II31694;
wire g12002;
wire II21494;
wire g24535;
wire II34274;
wire II40736;
wire g25421;
wire g27316;
wire g28045;
wire g24251;
wire II36981;
wire g13091;
wire g11652;
wire g21242;
wire g18379;
wire g5590;
wire II24694;
wire II23198;
wire g8178;
wire g9005;
wire II30302;
wire g5056;
wire II23605;
wire g16335;
wire g15424;
wire g10199;
wire g13411;
wire g29105;
wire II27164;
wire g5827;
wire II25831;
wire g7990;
wire g20728;
wire g25637;
wire II32424;
wire g23290;
wire II22902;
wire g29247;
wire g10497;
wire II15517;
wire g23495;
wire II23066;
wire g26767;
wire II16624;
wire g26751;
wire g19855;
wire g22286;
wire g8706;
wire g27290;
wire g23671;
wire g15868;
wire II23842;
wire g29173;
wire g17029;
wire II27369;
wire g10705;
wire g17462;
wire g26304;
wire g3494;
wire g16970;
wire g28916;
wire g8424;
wire g8432;
wire g13647;
wire g23774;
wire g24064;
wire g15991;
wire g17555;
wire g17131;
wire g26695;
wire II36758;
wire g7703;
wire g11035;
wire II36557;
wire g21183;
wire II39062;
wire g7582;
wire II22730;
wire II29159;
wire II31631;
wire g13552;
wire g26938;
wire II21955;
wire II33128;
wire g12935;
wire g16843;
wire g30644;
wire II23233;
wire g4142;
wire II31913;
wire g28346;
wire II14957;
wire g23783;
wire II26276;
wire g21738;
wire g28379;
wire g21773;
wire II39788;
wire II30335;
wire g17613;
wire II33593;
wire g26641;
wire g20609;
wire II20571;
wire g10035;
wire g23478;
wire g29240;
wire g11902;
wire II30245;
wire g4885;
wire II23575;
wire g21752;
wire g5187;
wire g28448;
wire g23878;
wire g27735;
wire II30953;
wire g17135;
wire g21868;
wire g29812;
wire g29095;
wire g29273;
wire II18148;
wire g7964;
wire g10511;
wire g18256;
wire g22515;
wire II29070;
wire II24514;
wire g21062;
wire g9588;
wire g8347;
wire g25148;
wire g30961;
wire g20600;
wire g25270;
wire g28842;
wire g29909;
wire II16479;
wire g19607;
wire II32646;
wire g22198;
wire g27186;
wire II25135;
wire II22631;
wire g20837;
wire g30702;
wire g29330;
wire g18919;
wire g30847;
wire g18926;
wire II33700;
wire g11504;
wire g15622;
wire gbuf57;
wire g19056;
wire II29429;
wire g26733;
wire g17175;
wire II26593;
wire II39779;
wire II38767;
wire g10323;
wire gbuf1;
wire g13944;
wire g24259;
wire II30948;
wire g8547;
wire g26043;
wire g20280;
wire g4313;
wire g6017;
wire g21861;
wire g23454;
wire II15369;
wire g4963;
wire II23661;
wire g10403;
wire g13991;
wire II15168;
wire g16292;
wire g26054;
wire II39323;
wire g22115;
wire g9010;
wire II24553;
wire g15971;
wire g18995;
wire g9368;
wire g30497;
wire g4705;
wire g15375;
wire g8135;
wire g20380;
wire g19905;
wire II24007;
wire g29031;
wire g28248;
wire II18271;
wire g30332;
wire g3937;
wire g13336;
wire g22264;
wire g17752;
wire g24735;
wire II31511;
wire g8528;
wire g29930;
wire II15015;
wire g28639;
wire g16102;
wire g23836;
wire g27331;
wire g13539;
wire II24016;
wire g22879;
wire g26779;
wire II30922;
wire g30814;
wire g22268;
wire g24012;
wire g14135;
wire II28975;
wire g13136;
wire g20944;
wire g13351;
wire g4775;
wire g12564;
wire g27416;
wire g19230;
wire g5770;
wire II14381;
wire II35067;
wire g13437;
wire II31036;
wire g26410;
wire g29146;
wire g19626;
wire g24563;
wire g7134;
wire g26772;
wire g16443;
wire g9723;
wire g26808;
wire g29782;
wire g10766;
wire g16791;
wire g28482;
wire g28241;
wire II17907;
wire II36577;
wire g5414;
wire g12128;
wire II18536;
wire g18646;
wire g25891;
wire g20590;
wire II34128;
wire g16478;
wire g24394;
wire g16462;
wire II29243;
wire II18494;
wire g18813;
wire g5919;
wire g17675;
wire g24825;
wire g18261;
wire g10492;
wire g28410;
wire g11768;
wire g11922;
wire g30057;
wire g21144;
wire g25593;
wire II14083;
wire g26714;
wire g13034;
wire g21782;
wire II40928;
wire g17713;
wire g30281;
wire II38160;
wire II25192;
wire II16549;
wire g10085;
wire g11877;
wire g10674;
wire g14963;
wire g28848;
wire g12966;
wire g27425;
wire g16438;
wire g24330;
wire g6103;
wire g12695;
wire g24633;
wire g14894;
wire g29311;
wire g30780;
wire g22710;
wire g30069;
wire g10952;
wire g4214;
wire g19401;
wire g19543;
wire II36237;
wire g28617;
wire g9047;
wire g29392;
wire g12211;
wire g10936;
wire II37858;
wire g18035;
wire g27293;
wire g9581;
wire g5297;
wire g27152;
wire g15781;
wire g9033;
wire g26271;
wire g24527;
wire g24266;
wire II23000;
wire g25565;
wire g16035;
wire g27082;
wire II13242;
wire g8939;
wire g17854;
wire g26687;
wire II23181;
wire g30207;
wire II36588;
wire g16284;
wire g15329;
wire g24363;
wire II20580;
wire g12866;
wire g28404;
wire II31571;
wire g18204;
wire II32528;
wire II18794;
wire g22316;
wire II31250;
wire g27385;
wire g27270;
wire g30346;
wire g26677;
wire g17988;
wire g26388;
wire g29636;
wire II39160;
wire g26665;
wire g23983;
wire g24908;
wire g15788;
wire g18332;
wire II38731;
wire g11815;
wire II25939;
wire II15787;
wire II29304;
wire g20739;
wire g7715;
wire g21564;
wire II20021;
wire g29797;
wire g23247;
wire g5104;
wire g11447;
wire g22680;
wire g11205;
wire g12448;
wire g21429;
wire g7748;
wire g17387;
wire g25038;
wire g5425;
wire II30914;
wire II33535;
wire g15685;
wire g26922;
wire II40856;
wire II16661;
wire II35900;
wire II32635;
wire g23387;
wire II16212;
wire g28154;
wire g9103;
wire II25846;
wire II35283;
wire II29206;
wire g23007;
wire II40853;
wire g19297;
wire g10614;
wire g28736;
wire g10292;
wire g9226;
wire g16775;
wire g25112;
wire g10209;
wire g29337;
wire g8871;
wire g16158;
wire g25935;
wire II18365;
wire g13406;
wire g27139;
wire II32880;
wire g26585;
wire g20990;
wire g21130;
wire g26481;
wire g5335;
wire g24958;
wire g30450;
wire II21392;
wire g30637;
wire II28491;
wire g15449;
wire II38885;
wire II19915;
wire g27037;
wire g15509;
wire g27447;
wire g7924;
wire II30782;
wire g27026;
wire II20685;
wire g9216;
wire II27516;
wire g4376;
wire g26998;
wire II34692;
wire g19295;
wire II34957;
wire II18665;
wire II17433;
wire II39878;
wire g27580;
wire g13278;
wire g28959;
wire g21761;
wire II28753;
wire g15055;
wire g12780;
wire II14541;
wire g22585;
wire g29367;
wire II33855;
wire g10862;
wire g23890;
wire II23976;
wire g27370;
wire g26288;
wire g30405;
wire g21634;
wire g8372;
wire g7922;
wire g28314;
wire g21529;
wire g22648;
wire g26630;
wire g24883;
wire g11858;
wire II37942;
wire g8816;
wire g22703;
wire g23098;
wire II38677;
wire g10202;
wire II16315;
wire g13871;
wire g21938;
wire g21096;
wire g5972;
wire g29046;
wire II31721;
wire II17151;
wire g30727;
wire g13213;
wire II26337;
wire g10422;
wire g19619;
wire g11674;
wire g4911;
wire g16662;
wire II16826;
wire II21884;
wire II32167;
wire II37415;
wire g12026;
wire g22812;
wire II19516;
wire g29201;
wire g17974;
wire g19187;
wire g10728;
wire g13067;
wire g11395;
wire II17831;
wire g13262;
wire g8825;
wire g5802;
wire II17012;
wire g4665;
wire g27507;
wire g15477;
wire g9528;
wire II25792;
wire g22043;
wire g8955;
wire II15267;
wire g23228;
wire g12542;
wire II24157;
wire II34438;
wire II36108;
wire g13180;
wire g25697;
wire g19112;
wire g30830;
wire g11748;
wire II40426;
wire g21392;
wire g20384;
wire g17307;
wire g30016;
wire g17094;
wire g11379;
wire g9118;
wire g29087;
wire g8182;
wire g8369;
wire g22954;
wire g10983;
wire II29129;
wire g21030;
wire g10390;
wire g12891;
wire II20505;
wire g27333;
wire g27030;
wire g30320;
wire II20394;
wire g30280;
wire g20560;
wire g22916;
wire g11129;
wire II21075;
wire II27727;
wire g26910;
wire g4721;
wire g10830;
wire g23510;
wire g24325;
wire g5645;
wire g19737;
wire II15278;
wire II33282;
wire g29630;
wire g30621;
wire g12961;
wire g24302;
wire g19368;
wire II18040;
wire g30856;
wire g28437;
wire g11608;
wire II31475;
wire g8482;
wire g15835;
wire II40438;
wire g19412;
wire g13050;
wire g26425;
wire g28987;
wire g26069;
wire g25963;
wire g26745;
wire g12192;
wire g26688;
wire g14016;
wire g4052;
wire g19247;
wire g29748;
wire g24518;
wire g13082;
wire g4073;
wire II30062;
wire II37467;
wire g7788;
wire g25991;
wire II34469;
wire g29289;
wire g5123;
wire g26205;
wire g5789;
wire g6517;
wire g23584;
wire g10271;
wire g19520;
wire II13652;
wire g8771;
wire II18704;
wire g22687;
wire g10073;
wire g19635;
wire g19173;
wire g27694;
wire II16736;
wire g27148;
wire g27286;
wire II17939;
wire g18424;
wire g29813;
wire II19836;
wire g18179;
wire g5902;
wire g10680;
wire g4092;
wire g11318;
wire II35796;
wire II31616;
wire g21042;
wire g21082;
wire g22400;
wire g30114;
wire g17186;
wire II16493;
wire g13636;
wire II33798;
wire g21671;
wire g5126;
wire g28423;
wire II14783;
wire II33891;
wire gbuf45;
wire II40895;
wire II39279;
wire II24279;
wire g13087;
wire g29224;
wire g30085;
wire g9077;
wire g8601;
wire g12555;
wire g21351;
wire g28648;
wire II24973;
wire g21047;
wire g4325;
wire g11987;
wire g23969;
wire g30679;
wire g5896;
wire II32490;
wire II26682;
wire g19949;
wire g20662;
wire g20597;
wire g29693;
wire g22662;
wire g29626;
wire II20538;
wire g19641;
wire g5153;
wire II34767;
wire II15237;
wire g5679;
wire II36797;
wire g12654;
wire g6711;
wire II14885;
wire g22911;
wire g26391;
wire II18079;
wire g12849;
wire g12382;
wire g23904;
wire g24830;
wire g27160;
wire g27130;
wire II31730;
wire II21432;
wire II22963;
wire g23688;
wire g17528;
wire g13448;
wire II21267;
wire g13106;
wire g5176;
wire g28419;
wire g21358;
wire g5834;
wire II24374;
wire g18070;
wire g27103;
wire gbuf38;
wire g28464;
wire II16012;
wire II29162;
wire g14008;
wire g23661;
wire g25251;
wire g30907;
wire II15605;
wire g27886;
wire g20331;
wire II15559;
wire g10435;
wire II23124;
wire II21601;
wire g4243;
wire g29513;
wire II38743;
wire II23094;
wire g8458;
wire g21449;
wire g16852;
wire g28283;
wire g5658;
wire II18408;
wire g13365;
wire g26596;
wire II18073;
wire II27011;
wire g24029;
wire II29010;
wire g26955;
wire g15731;
wire g9711;
wire g18605;
wire II28031;
wire II38647;
wire g22075;
wire g7900;
wire II21705;
wire gbuf40;
wire g10443;
wire g10904;
wire II32857;
wire g20613;
wire II22926;
wire II28217;
wire g24409;
wire II30676;
wire g28027;
wire g12882;
wire II34135;
wire II22771;
wire II22539;
wire g23694;
wire g13129;
wire g28432;
wire gbuf29;
wire g22218;
wire II23851;
wire II24195;
wire II40300;
wire g21659;
wire g4728;
wire g9757;
wire g13918;
wire g29790;
wire g25479;
wire g30808;
wire II38505;
wire g15738;
wire g20874;
wire g18311;
wire g29767;
wire g12170;
wire g28525;
wire g24575;
wire g15959;
wire g27171;
wire g8200;
wire g19702;
wire g26662;
wire g28322;
wire II35431;
wire gbuf22;
wire g23279;
wire g4121;
wire g10360;
wire g30944;
wire g5469;
wire g19809;
wire g28071;
wire g11889;
wire II23383;
wire g17402;
wire II31008;
wire g28104;
wire g19804;
wire g7629;
wire g14062;
wire II40537;
wire II35172;
wire g21022;
wire II39475;
wire g8099;
wire g5761;
wire g16865;
wire II18386;
wire II18644;
wire g5720;
wire g16988;
wire g28392;
wire II25572;
wire g27502;
wire g13674;
wire g8553;
wire g18945;
wire g14881;
wire g20313;
wire g26220;
wire g17247;
wire g30698;
wire II18061;
wire g22151;
wire g14165;
wire g6369;
wire g23729;
wire g28376;
wire g30372;
wire g22166;
wire II29026;
wire g26982;
wire g29424;
wire II19820;
wire g13170;
wire g28725;
wire g21002;
wire g21875;
wire g18856;
wire g5401;
wire g13862;
wire II19315;
wire g6978;
wire g19158;
wire g21079;
wire g26823;
wire g18504;
wire II37760;
wire II16650;
wire g12790;
wire g23919;
wire g15550;
wire g28062;
wire II34369;
wire g29466;
wire g19233;
wire g10901;
wire II25811;
wire g15196;
wire g15923;
wire g12426;
wire g17566;
wire g13568;
wire g14442;
wire g28762;
wire g10389;
wire g20156;
wire g17142;
wire g29487;
wire g28584;
wire II14819;
wire g16177;
wire g28005;
wire g7812;
wire g7827;
wire II35879;
wire II29191;
wire g19021;
wire g30248;
wire g11498;
wire g16040;
wire II25399;
wire g24648;
wire g11717;
wire g29433;
wire g24335;
wire g19595;
wire g26604;
wire II20425;
wire g22832;
wire g12950;
wire g27823;
wire g26883;
wire II20117;
wire g23242;
wire g9507;
wire g12264;
wire g10047;
wire II15584;
wire g6943;
wire g20438;
wire g26426;
wire II36502;
wire II36891;
wire g26446;
wire g8027;
wire g17240;
wire g19151;
wire g9050;
wire II23521;
wire g24820;
wire II22836;
wire g19838;
wire g20360;
wire g27514;
wire g19093;
wire g28353;
wire g9425;
wire g23050;
wire g26884;
wire g13699;
wire g29769;
wire g4753;
wire II30152;
wire g19864;
wire g27533;
wire g12177;
wire II40456;
wire g18622;
wire g7822;
wire II26541;
wire g19494;
wire g16415;
wire g19279;
wire g27703;
wire g12822;
wire g19742;
wire g30363;
wire g13859;
wire g24067;
wire g30354;
wire g8083;
wire g29475;
wire g29972;
wire II30050;
wire II39133;
wire g3410;
wire g11566;
wire g24056;
wire g10185;
wire g24486;
wire g15337;
wire II29562;
wire g25033;
wire II37897;
wire g19929;
wire g15525;
wire g24586;
wire g26192;
wire g13511;
wire g24492;
wire g28253;
wire g6220;
wire g30125;
wire g25968;
wire gbuf182;
wire g23216;
wire g24520;
wire g28399;
wire g13962;
wire g25059;
wire g28729;
wire g26504;
wire g21203;
wire g15126;
wire II33861;
wire II17948;
wire g12596;
wire II25607;
wire g11675;
wire II36090;
wire g27797;
wire g20410;
wire g26891;
wire g11824;
wire II21108;
wire g24857;
wire g26489;
wire g7760;
wire g12220;
wire g21483;
wire g21308;
wire g25395;
wire g4587;
wire g9260;
wire II28981;
wire g30467;
wire g16065;
wire II23599;
wire g6284;
wire II15568;
wire II23490;
wire g9884;
wire g12457;
wire g16412;
wire II40754;
wire g13159;
wire g26125;
wire g24448;
wire g13756;
wire g26348;
wire g15792;
wire g19253;
wire II40742;
wire g26020;
wire g14408;
wire g15248;
wire g27632;
wire g19269;
wire g19193;
wire II28512;
wire g20810;
wire g9504;
wire g4620;
wire g12218;
wire g29917;
wire g19760;
wire g30762;
wire g21168;
wire II21666;
wire g15698;
wire g27253;
wire g26989;
wire II22584;
wire g30266;
wire g10282;
wire g11832;
wire g10119;
wire g16429;
wire g26150;
wire g23274;
wire g24471;
wire gbuf178;
wire g22387;
wire g13295;
wire g21892;
wire g24236;
wire g18963;
wire g8062;
wire g30100;
wire g15729;
wire g26873;
wire g13044;
wire g20980;
wire II34641;
wire g22228;
wire g16475;
wire II32949;
wire g10835;
wire g20687;
wire g19881;
wire II14295;
wire g15343;
wire g29670;
wire g10637;
wire g30454;
wire g30672;
wire II40763;
wire g16659;
wire g28670;
wire g26974;
wire g27770;
wire g12166;
wire g13990;
wire g27542;
wire g19260;
wire g15813;
wire g29290;
wire g16223;
wire g22029;
wire g19652;
wire g19822;
wire g8687;
wire g21444;
wire g29157;
wire II35762;
wire g17544;
wire g16419;
wire II20295;
wire g25088;
wire II27122;
wire g26543;
wire g5024;
wire II16514;
wire g25524;
wire g21266;
wire g16075;
wire g7892;
wire II21739;
wire g25130;
wire g20316;
wire g28686;
wire II33437;
wire g23065;
wire II36397;
wire g3951;
wire II15810;
wire g30650;
wire g29910;
wire g8447;
wire g21445;
wire g21968;
wire g21267;
wire g25672;
wire g18240;
wire II20616;
wire g19217;
wire II23095;
wire g30657;
wire g24459;
wire g8191;
wire II31892;
wire g19038;
wire g28268;
wire II33912;
wire II24252;
wire g30683;
wire II37746;
wire g19757;
wire gbuf105;
wire g28189;
wire g30077;
wire g27118;
wire g24450;
wire g20019;
wire II32085;
wire g29268;
wire g15780;
wire g19186;
wire II20355;
wire g11673;
wire g20198;
wire II29954;
wire II21962;
wire II31559;
wire g28009;
wire g24090;
wire II31469;
wire g9569;
wire gbuf93;
wire g20995;
wire g29897;
wire g5729;
wire II17184;
wire gbuf117;
wire g15326;
wire II18396;
wire g17324;
wire g28634;
wire g23687;
wire g24760;
wire II37851;
wire g28243;
wire g12441;
wire g27766;
wire II14163;
wire g16277;
wire g7911;
wire g6201;
wire g5925;
wire g14507;
wire II27832;
wire II21326;
wire g26400;
wire II31844;
wire g30017;
wire g10585;
wire g11092;
wire g29010;
wire g11845;
wire g11879;
wire g26373;
wire g13815;
wire II27246;
wire g15787;
wire g15641;
wire g20894;
wire g27497;
wire g18821;
wire g4623;
wire g19251;
wire II25635;
wire II36315;
wire g5680;
wire g4197;
wire II32617;
wire g13825;
wire g3554;
wire g12993;
wire g15842;
wire g8892;
wire II37311;
wire g23251;
wire II13207;
wire g24815;
wire g4009;
wire g3366;
wire g24264;
wire g18941;
wire g16360;
wire II19898;
wire II18308;
wire g10174;
wire g29582;
wire g12242;
wire g29107;
wire g28372;
wire g5765;
wire g18830;
wire g27526;
wire g15811;
wire g5874;
wire gbuf75;
wire g21189;
wire g15106;
wire g19248;
wire g24222;
wire g28396;
wire g14669;
wire g20293;
wire g11681;
wire g20973;
wire g4956;
wire gbuf179;
wire II21758;
wire g24791;
wire II21297;
wire g14297;
wire II26266;
wire g28694;
wire g17022;
wire g29982;
wire g27383;
wire II27976;
wire g23348;
wire II33312;
wire II34266;
wire II31760;
wire g29834;
wire g8780;
wire II31796;
wire g22148;
wire g30520;
wire g30513;
wire g21750;
wire g18401;
wire g26438;
wire g13032;
wire II37173;
wire g4091;
wire II36679;
wire g12065;
wire g5983;
wire g29817;
wire II19513;
wire II32281;
wire g13294;
wire g13884;
wire g11942;
wire g19166;
wire II22936;
wire II33834;
wire II27614;
wire g13526;
wire II15205;
wire g10681;
wire g21276;
wire II25605;
wire g20134;
wire g20601;
wire II29226;
wire II31652;
wire g8075;
wire g24338;
wire II19816;
wire II20679;
wire g14061;
wire g25923;
wire II26420;
wire g13126;
wire g25149;
wire g29495;
wire g24776;
wire g10784;
wire g11722;
wire g30699;
wire g30583;
wire g25004;
wire g13248;
wire g6942;
wire g30730;
wire II18770;
wire g19199;
wire g28784;
wire g9767;
wire g23306;
wire g27999;
wire g8385;
wire g23088;
wire II25654;
wire II16641;
wire II23314;
wire II30888;
wire g26769;
wire g17619;
wire g26999;
wire II24646;
wire g21882;
wire g23453;
wire g12216;
wire g4526;
wire g16130;
wire g7158;
wire g8757;
wire g30062;
wire g30007;
wire g12196;
wire g22551;
wire g16238;
wire g21285;
wire g26849;
wire II23358;
wire g22833;
wire II16267;
wire II22964;
wire g11595;
wire II29588;
wire II20031;
wire g25648;
wire II16578;
wire g28128;
wire II34845;
wire g18638;
wire g28354;
wire g4644;
wire g19857;
wire II35667;
wire II15475;
wire g13724;
wire g28471;
wire g24099;
wire g23195;
wire g23795;
wire II19274;
wire II24612;
wire II38477;
wire g25023;
wire g25066;
wire g11514;
wire g14412;
wire II13200;
wire II14665;
wire g25180;
wire II26621;
wire g15826;
wire g26000;
wire g4839;
wire g18448;
wire g18030;
wire g4208;
wire g20517;
wire g26534;
wire II22560;
wire g13076;
wire g26621;
wire II32895;
wire g22434;
wire g25365;
wire II19767;
wire g21031;
wire g7936;
wire II25681;
wire g20676;
wire g21057;
wire g16636;
wire g17557;
wire g19078;
wire II31643;
wire g28017;
wire II28458;
wire g11507;
wire g26752;
wire g10606;
wire g22013;
wire g20054;
wire g29521;
wire g18585;
wire g28086;
wire g17508;
wire g12534;
wire g19387;
wire g13355;
wire g19080;
wire g16471;
wire II39341;
wire g28103;
wire g27094;
wire g20628;
wire II14650;
wire II24091;
wire g20312;
wire g21258;
wire II33355;
wire II32175;
wire g14650;
wire g5141;
wire g22880;
wire g18142;
wire II25673;
wire g14206;
wire g30044;
wire II40685;
wire g16123;
wire g5269;
wire g8766;
wire g6065;
wire g21957;
wire g16862;
wire II24487;
wire g22291;
wire II23611;
wire II29119;
wire gbuf46;
wire g28320;
wire g28527;
wire g20327;
wire II16782;
wire g26628;
wire g14493;
wire g15505;
wire g11993;
wire g30960;
wire II25723;
wire II14553;
wire g12290;
wire g10963;
wire g7539;
wire II18353;
wire g30927;
wire g4603;
wire II41102;
wire II40558;
wire II36792;
wire g26392;
wire g30839;
wire g15488;
wire g27162;
wire II29277;
wire g30853;
wire II16050;
wire g22704;
wire g30310;
wire II17712;
wire g27366;
wire g25312;
wire g11401;
wire g17348;
wire g12055;
wire g19669;
wire g30610;
wire g12989;
wire g5047;
wire g20565;
wire g30025;
wire g10286;
wire II25492;
wire II28111;
wire g24462;
wire g22030;
wire g30319;
wire g30969;
wire g12408;
wire II30511;
wire g24297;
wire g25953;
wire g25252;
wire g21372;
wire g5916;
wire g29780;
wire II28191;
wire g16817;
wire g23423;
wire II34788;
wire g19027;
wire g22057;
wire II34056;
wire II26388;
wire g19677;
wire g15855;
wire g22025;
wire II40868;
wire II24711;
wire g19673;
wire g26172;
wire g21813;
wire g21071;
wire II38355;
wire g4803;
wire g24107;
wire g19328;
wire g18153;
wire g26563;
wire g11620;
wire g27765;
wire g8324;
wire g28484;
wire g27278;
wire g9872;
wire g21920;
wire II14580;
wire g19670;
wire g17160;
wire II38609;
wire g8045;
wire II19479;
wire II29972;
wire g29414;
wire g9203;
wire g11833;
wire g28700;
wire g22437;
wire g18869;
wire g20935;
wire g19534;
wire g22720;
wire g15390;
wire g3772;
wire II30167;
wire g18047;
wire g24537;
wire g24082;
wire g22665;
wire II29110;
wire g24100;
wire g25746;
wire g23269;
wire g11014;
wire g9093;
wire g10516;
wire g27051;
wire g30805;
wire g23206;
wire II17813;
wire g17990;
wire g11558;
wire g14467;
wire II39411;
wire g4029;
wire g18484;
wire g24731;
wire g25643;
wire g30124;
wire g25341;
wire II30035;
wire II26972;
wire g20353;
wire g29507;
wire g29035;
wire g3834;
wire g21927;
wire g20161;
wire II18479;
wire II16936;
wire g30370;
wire g21331;
wire g9122;
wire g5601;
wire g5548;
wire II17843;
wire g23769;
wire II37484;
wire II13137;
wire II34653;
wire g23511;
wire II30275;
wire g30782;
wire g28118;
wire II22019;
wire g4012;
wire g30860;
wire g21851;
wire II23190;
wire g19205;
wire g24595;
wire g17327;
wire g30936;
wire g5948;
wire g15188;
wire g16633;
wire g18542;
wire g30822;
wire g13476;
wire g23895;
wire g27869;
wire II18326;
wire II32925;
wire g18873;
wire g24133;
wire g11854;
wire g28047;
wire g8168;
wire g13613;
wire g13374;
wire g13895;
wire g9232;
wire g27218;
wire g10309;
wire g27058;
wire g9084;
wire g16989;
wire g29527;
wire g17696;
wire g24861;
wire II23398;
wire g6301;
wire g5996;
wire g29061;
wire g10831;
wire g6197;
wire g26598;
wire g11389;
wire II27385;
wire II16897;
wire g20038;
wire II25616;
wire g30617;
wire g23104;
wire g29702;
wire g7328;
wire g8302;
wire II38728;
wire g17648;
wire g17235;
wire g7424;
wire g16097;
wire g19568;
wire g17390;
wire II26240;
wire g9319;
wire g26103;
wire II34444;
wire II24657;
wire g12601;
wire g8246;
wire g29731;
wire II27152;
wire g24986;
wire II30792;
wire g29085;
wire g11962;
wire II38111;
wire II22587;
wire g22811;
wire II23542;
wire g22167;
wire g22718;
wire g5333;
wire g9926;
wire II21780;
wire g22404;
wire II36227;
wire g25874;
wire g10017;
wire g24541;
wire II24465;
wire g10416;
wire g4188;
wire g13268;
wire g13836;
wire II21395;
wire g28657;
wire g28254;
wire g8245;
wire g11892;
wire g22550;
wire g5421;
wire g19893;
wire II40880;
wire g23664;
wire g19019;
wire g12030;
wire g17230;
wire g29779;
wire g25691;
wire g16495;
wire g22646;
wire g18497;
wire II19595;
wire g13852;
wire g27229;
wire II18414;
wire g16823;
wire g12828;
wire g24123;
wire g14702;
wire g17610;
wire II38764;
wire g29617;
wire II36684;
wire g10146;
wire g29335;
wire g25467;
wire II13146;
wire g26824;
wire II18800;
wire g27359;
wire g13066;
wire g20405;
wire g4595;
wire II14634;
wire g9480;
wire II27372;
wire g20426;
wire g3966;
wire II16879;
wire g23580;
wire g27950;
wire g13739;
wire g22632;
wire g16348;
wire g6444;
wire II14513;
wire II29516;
wire II30323;
wire g19477;
wire g15350;
wire g19875;
wire g27919;
wire g26246;
wire g22464;
wire II24738;
wire g5004;
wire g22365;
wire II23633;
wire II18088;
wire g5797;
wire g19698;
wire g29089;
wire g28719;
wire g26602;
wire g10474;
wire g18514;
wire g24878;
wire g7162;
wire g30018;
wire II33368;
wire g20184;
wire g24545;
wire g23096;
wire II40002;
wire g4061;
wire II23782;
wire II29663;
wire II17792;
wire g27882;
wire II40700;
wire g22850;
wire g26488;
wire II38629;
wire II22982;
wire g24851;
wire II20410;
wire II23104;
wire g8823;
wire g12971;
wire II15244;
wire g30976;
wire II40581;
wire g30290;
wire g29532;
wire g18665;
wire II19808;
wire g22239;
wire II16966;
wire g5358;
wire g15547;
wire g5855;
wire g11773;
wire g24840;
wire g27001;
wire II40248;
wire g28553;
wire g10871;
wire g26890;
wire g27712;
wire g10467;
wire II40027;
wire II14842;
wire II38770;
wire g12274;
wire g19885;
wire II32129;
wire g16058;
wire g8578;
wire g22298;
wire II30347;
wire II35509;
wire g26292;
wire g15777;
wire g17297;
wire g9603;
wire g18937;
wire II28541;
wire g26021;
wire g26685;
wire g22037;
wire g23364;
wire g27928;
wire II14981;
wire g30834;
wire II37924;
wire II22515;
wire II32510;
wire II31514;
wire g26164;
wire II35837;
wire g11564;
wire g23071;
wire II18338;
wire g18643;
wire g15052;
wire g10851;
wire II36129;
wire g24051;
wire g13657;
wire g25105;
wire g14454;
wire g28924;
wire II25486;
wire g11471;
wire II21878;
wire II38843;
wire II27047;
wire g23838;
wire g27509;
wire g16388;
wire g12439;
wire g22315;
wire g30031;
wire II27288;
wire II32527;
wire g28369;
wire g15271;
wire II31610;
wire II34327;
wire g27261;
wire g9636;
wire g25612;
wire g24410;
wire g27686;
wire II24103;
wire g24350;
wire g25318;
wire g20574;
wire g28662;
wire g11546;
wire g27801;
wire II28467;
wire g29419;
wire g27282;
wire g8144;
wire II38638;
wire g16467;
wire g8516;
wire g29718;
wire g19572;
wire g22170;
wire g21134;
wire g5009;
wire g24564;
wire g16832;
wire II14472;
wire g9961;
wire g25771;
wire g8972;
wire g5319;
wire g9940;
wire g11111;
wire II20520;
wire g26720;
wire g28409;
wire g23184;
wire II33846;
wire g3972;
wire II35983;
wire II27086;
wire g19325;
wire g28833;
wire g19519;
wire II25866;
wire II18191;
wire g12867;
wire g29429;
wire g8507;
wire g28037;
wire II37653;
wire g18355;
wire g9354;
wire g9245;
wire g10929;
wire II37080;
wire g5967;
wire g22788;
wire g22226;
wire g30111;
wire g21199;
wire II32688;
wire g6135;
wire g20666;
wire II36879;
wire II20050;
wire g13970;
wire g14956;
wire g8580;
wire g13291;
wire II35072;
wire g30796;
wire g30483;
wire II19727;
wire II30589;
wire g22339;
wire II38042;
wire g4156;
wire g17813;
wire g7556;
wire g9622;
wire g26541;
wire g11144;
wire g13643;
wire II28742;
wire g9035;
wire g25262;
wire g11521;
wire II32538;
wire II19637;
wire II17641;
wire g11817;
wire g7606;
wire g21931;
wire g6427;
wire g13459;
wire II34921;
wire g23029;
wire g24494;
wire g16199;
wire g10694;
wire II29490;
wire g12151;
wire II30496;
wire g24839;
wire g24395;
wire g15171;
wire g9902;
wire II28013;
wire g10482;
wire g27450;
wire g14395;
wire g21486;
wire g27070;
wire g15581;
wire g29929;
wire g14113;
wire II25821;
wire II26220;
wire g6896;
wire II16984;
wire g29649;
wire g26099;
wire II29432;
wire g28397;
wire II32324;
wire g24929;
wire g7757;
wire g13672;
wire II25539;
wire g23060;
wire g18447;
wire II33418;
wire g8469;
wire II31532;
wire g26868;
wire g11790;
wire g26729;
wire g24912;
wire II31925;
wire g26339;
wire g24206;
wire g22344;
wire g12178;
wire g30446;
wire II18838;
wire II30242;
wire g11806;
wire g30303;
wire g10311;
wire g15721;
wire g23521;
wire g29030;
wire g8863;
wire g24361;
wire II40504;
wire g29212;
wire II18253;
wire g10133;
wire II25865;
wire II31235;
wire II37778;
wire g26046;
wire g9465;
wire II34974;
wire g10660;
wire g26804;
wire g27206;
wire g4898;
wire g21966;
wire g12642;
wire g8940;
wire g7149;
wire g13461;
wire g27155;
wire g16999;
wire II35011;
wire II37089;
wire g19622;
wire g28343;
wire g17129;
wire g22087;
wire g13588;
wire g16854;
wire g23502;
wire g25115;
wire g30330;
wire g20918;
wire II25596;
wire g30492;
wire II40697;
wire g13137;
wire g8239;
wire g9629;
wire g16990;
wire g23486;
wire g25322;
wire II15827;
wire g21576;
wire g30815;
wire g15719;
wire g21233;
wire g26449;
wire g27660;
wire g25862;
wire II41041;
wire II36490;
wire g8164;
wire II33567;
wire II29148;
wire II15451;
wire II24704;
wire g13313;
wire g18822;
wire g29174;
wire g11732;
wire g12185;
wire g5289;
wire II38686;
wire g22840;
wire g29822;
wire g17363;
wire g19545;
wire g30827;
wire g23440;
wire g5610;
wire g26036;
wire II17762;
wire g23527;
wire g9610;
wire g27106;
wire g17868;
wire g12377;
wire g28608;
wire g10037;
wire II15925;
wire g11952;
wire g27532;
wire g11617;
wire II30832;
wire II36554;
wire g12049;
wire g20535;
wire g28030;
wire g11154;
wire II20661;
wire g23537;
wire g4778;
wire II38665;
wire g26780;
wire g5372;
wire g19915;
wire II25665;
wire g23296;
wire g21052;
wire g28028;
wire g3963;
wire g30437;
wire g11851;
wire g16067;
wire g26827;
wire II21641;
wire g26092;
wire g11585;
wire g30345;
wire II17740;
wire g21658;
wire II23409;
wire g8437;
wire g17598;
wire g16139;
wire g16073;
wire g5974;
wire g29150;
wire g26833;
wire II37813;
wire g18333;
wire g24956;
wire g8025;
wire g6363;
wire II15487;
wire g15872;
wire g22076;
wire g29443;
wire II27303;
wire II38097;
wire g23444;
wire g29962;
wire g24795;
wire II28076;
wire II29402;
wire II40518;
wire g6035;
wire g18785;
wire g19601;
wire g26131;
wire g7595;
wire g17838;
wire g30257;
wire II16354;
wire II35059;
wire g20881;
wire II29993;
wire g23142;
wire II28833;
wire g15707;
wire g19102;
wire g13561;
wire g30395;
wire g26805;
wire g19715;
wire II36483;
wire g14144;
wire g7796;
wire g11574;
wire II40844;
wire g12171;
wire g5943;
wire g17220;
wire g15901;
wire g8534;
wire g12308;
wire g21877;
wire g26361;
wire g16219;
wire g30360;
wire II35057;
wire II19530;
wire g27847;
wire g21945;
wire g10793;
wire g17600;
wire g16163;
wire g6156;
wire g6141;
wire II38077;
wire II19380;
wire II26714;
wire g30947;
wire II33466;
wire g18388;
wire g12331;
wire II18767;
wire g30571;
wire II30816;
wire g17176;
wire II34183;
wire g11698;
wire g19561;
wire g26676;
wire g27211;
wire g27285;
wire g25811;
wire g7615;
wire g5709;
wire g7592;
wire g22195;
wire g21015;
wire g23634;
wire g22443;
wire g10273;
wire II16079;
wire g4047;
wire g29258;
wire g30881;
wire II30686;
wire g11456;
wire II32901;
wire II40823;
wire g12598;
wire g29233;
wire g20272;
wire g28236;
wire g29210;
wire g29287;
wire g22772;
wire g30848;
wire g19860;
wire g5863;
wire g7971;
wire g6678;
wire g28388;
wire g14472;
wire g15763;
wire g19608;
wire g28495;
wire g26914;
wire g25661;
wire II41120;
wire g12967;
wire g21305;
wire g8905;
wire g8630;
wire g17962;
wire g29640;
wire g28951;
wire II25246;
wire II21482;
wire II30116;
wire g22230;
wire g25626;
wire g29942;
wire g23578;
wire II28443;
wire g11821;
wire g28302;
wire g20672;
wire g22255;
wire g10383;
wire II30707;
wire g22670;
wire g23739;
wire g28723;
wire g16743;
wire g18885;
wire II32647;
wire g6572;
wire g9009;
wire g15228;
wire g30778;
wire g8277;
wire g27436;
wire g17158;
wire g30757;
wire g25976;
wire g13021;
wire II32388;
wire II18121;
wire g29804;
wire g24599;
wire II23539;
wire g24616;
wire g24150;
wire g11939;
wire II29635;
wire g15287;
wire II18389;
wire g25993;
wire g19143;
wire g25164;
wire g22201;
wire g18464;
wire II22901;
wire g30246;
wire g24275;
wire g20375;
wire g23282;
wire II17721;
wire II16363;
wire g23940;
wire g23616;
wire g29566;
wire g16447;
wire II31027;
wire g10528;
wire II18268;
wire g8925;
wire g13869;
wire II33476;
wire g10197;
wire II41017;
wire II31062;
wire II25977;
wire II37702;
wire g8845;
wire g17123;
wire g20370;
wire g21907;
wire g22624;
wire g20000;
wire g6117;
wire II16312;
wire g30987;
wire g17984;
wire II41010;
wire g16381;
wire g16622;
wire g20945;
wire g13483;
wire II23045;
wire g27132;
wire g17902;
wire g19413;
wire II18671;
wire g25197;
wire g7733;
wire g27192;
wire g25452;
wire g13506;
wire g25061;
wire II31712;
wire g21111;
wire II27253;
wire g28478;
wire g27554;
wire g19305;
wire g5821;
wire g21177;
wire g13367;
wire g20591;
wire g19400;
wire g21900;
wire II28953;
wire g17966;
wire g13270;
wire II28500;
wire g26696;
wire g17487;
wire II32498;
wire g23916;
wire g28200;
wire II23857;
wire g25668;
wire g5196;
wire g6085;
wire g12565;
wire g12854;
wire g22448;
wire g27348;
wire II41066;
wire g19790;
wire g12156;
wire II18094;
wire g7849;
wire g21394;
wire g9382;
wire g28191;
wire g24805;
wire g21496;
wire gbuf107;
wire g20478;
wire g30592;
wire g5218;
wire g29310;
wire g6028;
wire g15941;
wire II35440;
wire II16633;
wire II29736;
wire g27916;
wire g30891;
wire g15502;
wire g17475;
wire g29954;
wire g21192;
wire g21980;
wire g29207;
wire II25532;
wire II24625;
wire II31257;
wire g5075;
wire II37098;
wire g25296;
wire g18597;
wire II32586;
wire g27074;
wire g7655;
wire g6173;
wire g10126;
wire g18846;
wire g18573;
wire g9531;
wire gbuf2;
wire g22251;
wire g23076;
wire g30439;
wire g18436;
wire g10508;
wire g22050;
wire II39764;
wire gbuf184;
wire g5883;
wire g12688;
wire g30799;
wire g22116;
wire g27924;
wire g27173;
wire g30560;
wire II39889;
wire g28040;
wire g26270;
wire II22569;
wire g11970;
wire g13849;
wire g23614;
wire g10779;
wire II34901;
wire g9049;
wire g13004;
wire g27965;
wire g30514;
wire g29662;
wire g10454;
wire II23602;
wire II37305;
wire g24419;
wire g27629;
wire g10462;
wire g11300;
wire II18602;
wire g23596;
wire g10062;
wire II33377;
wire g24847;
wire II20799;
wire g28454;
wire g30256;
wire II25064;
wire II18467;
wire g29479;
wire g30271;
wire g27945;
wire II29660;
wire g20954;
wire g13211;
wire g10537;
wire g22677;
wire g22042;
wire g18907;
wire II23019;
wire g13926;
wire g22415;
wire g29077;
wire g27576;
wire II29519;
wire g27245;
wire II23967;
wire g27302;
wire g20580;
wire II18668;
wire II39246;
wire II38827;
wire II21736;
wire g22795;
wire II31592;
wire II23010;
wire g19481;
wire g12949;
wire g23114;
wire g19775;
wire g13203;
wire g16092;
wire g29377;
wire g27409;
wire g20149;
wire II17103;
wire II20466;
wire g7455;
wire g10153;
wire II16244;
wire g7868;
wire g28109;
wire II40841;
wire II35389;
wire g26238;
wire g13114;
wire g23801;
wire g26356;
wire II40871;
wire g29359;
wire g26265;
wire g10530;
wire g30252;
wire g23546;
wire g29997;
wire g11670;
wire II33307;
wire II20278;
wire II35449;
wire g26212;
wire g11422;
wire g10912;
wire II16723;
wire II27179;
wire II33300;
wire g20044;
wire g23175;
wire g15418;
wire g19013;
wire g19977;
wire g28067;
wire II22699;
wire g11885;
wire g28384;
wire g10582;
wire g19616;
wire g26343;
wire II34009;
wire II39840;
wire g7975;
wire II40066;
wire II18539;
wire II34731;
wire g10908;
wire g12930;
wire g22138;
wire II25315;
wire g4363;
wire g10557;
wire g10376;
wire g29435;
wire g16242;
wire g29516;
wire g13284;
wire g15379;
wire II30200;
wire g20618;
wire g21971;
wire g26928;
wire g20749;
wire II23244;
wire II39976;
wire II38671;
wire g18976;
wire g27505;
wire g22279;
wire g13513;
wire g25919;
wire g28444;
wire g21043;
wire g4412;
wire g5752;
wire g22827;
wire g25707;
wire II36117;
wire II30293;
wire g28325;
wire II14584;
wire g27220;
wire II36966;
wire II21514;
wire g20158;
wire g23853;
wire g22455;
wire g20465;
wire g29497;
wire g22243;
wire gbuf100;
wire g22765;
wire g15402;
wire g21976;
wire g8977;
wire II27197;
wire g28004;
wire g8882;
wire II18656;
wire g30545;
wire g20191;
wire II38916;
wire g15833;
wire g5696;
wire g27698;
wire g19154;
wire g19090;
wire II31050;
wire g16213;
wire g9673;
wire g26931;
wire g26918;
wire II22823;
wire g19179;
wire g27691;
wire g30877;
wire g10905;
wire II18813;
wire g26786;
wire g30640;
wire II37620;
wire g15849;
wire g30447;
wire g20393;
wire g22636;
wire g20729;
wire g27550;
wire g14537;
wire g20277;
wire II22317;
wire II36766;
wire II19318;
wire II31880;
wire g13090;
wire II35876;
wire g12470;
wire gbuf205;
wire g19694;
wire g10593;
wire II16521;
wire g22124;
wire II20658;
wire g29461;
wire g30535;
wire g20912;
wire g7078;
wire g12175;
wire g17302;
wire g29741;
wire g21454;
wire g4246;
wire g27257;
wire II37875;
wire g27125;
wire g10747;
wire g20159;
wire II21655;
wire g14601;
wire g22155;
wire II39550;
wire g24166;
wire g13840;
wire II19545;
wire g10364;
wire II39267;
wire g9061;
wire g23685;
wire g7679;
wire g26836;
wire g29482;
wire II22707;
wire II33198;
wire II16144;
wire g7347;
wire g26042;
wire g12045;
wire g14849;
wire II24227;
wire g18522;
wire II26481;
wire II40682;
wire g13323;
wire g6183;
wire II32120;
wire g24653;
wire g30957;
wire II31871;
wire II39472;
wire II29405;
wire g19031;
wire II34192;
wire g12544;
wire g29463;
wire g18982;
wire g10858;
wire g27700;
wire g19547;
wire II21119;
wire II38369;
wire g11332;
wire g24232;
wire g27114;
wire g11801;
wire g5713;
wire g22612;
wire g30028;
wire g4292;
wire g3928;
wire g28737;
wire g17621;
wire g21202;
wire II31102;
wire g27830;
wire g18217;
wire g10627;
wire II25521;
wire g22570;
wire g18508;
wire g12453;
wire II24595;
wire II34041;
wire g11789;
wire II23518;
wire g16411;
wire g17413;
wire g29633;
wire g15921;
wire g11926;
wire g25037;
wire g5309;
wire g20742;
wire g12702;
wire II30029;
wire g28696;
wire g20434;
wire g19807;
wire g14040;
wire g19229;
wire II31634;
wire g28297;
wire g23594;
wire II36864;
wire g14768;
wire g20334;
wire g29294;
wire g30518;
wire g20587;
wire II23179;
wire g15724;
wire g13796;
wire g15325;
wire g8899;
wire g18853;
wire II28043;
wire g25399;
wire g4340;
wire II38142;
wire g28258;
wire g13936;
wire g10193;
wire g28810;
wire gbuf172;
wire g24886;
wire g24246;
wire g12490;
wire g21008;
wire g21480;
wire II19958;
wire g7138;
wire g17083;
wire g20997;
wire g23164;
wire g21209;
wire II30607;
wire g10361;
wire g15340;
wire g25964;
wire II40721;
wire g21987;
wire II17228;
wire g29279;
wire g19896;
wire g10829;
wire gbuf73;
wire g23110;
wire II40766;
wire II31478;
wire g13515;
wire g11661;
wire g23710;
wire g10122;
wire g28880;
wire II24180;
wire g10189;
wire g29613;
wire g26121;
wire II25712;
wire g21806;
wire g4329;
wire II37140;
wire g28075;
wire g17213;
wire II36733;
wire g18725;
wire g7897;
wire g20415;
wire g30932;
wire II33608;
wire g5327;
wire II25081;
wire g18244;
wire g28663;
wire g29885;
wire II24586;
wire g13153;
wire II30536;
wire II24668;
wire g4832;
wire II21775;
wire II15329;
wire II35515;
wire II20810;
wire g25134;
wire II27128;
wire g16152;
wire g21716;
wire II39407;
wire g16312;
wire g13039;
wire g21674;
wire g24578;
wire II23807;
wire II38499;
wire g8874;
wire g12900;
wire g26461;
wire g30359;
wire g13850;
wire II33013;
wire II35937;
wire g26996;
wire g26495;
wire g26775;
wire g24262;
wire g9400;
wire g12147;
wire g15846;
wire g27517;
wire g11982;
wire g13433;
wire g21847;
wire g26119;
wire g25549;
wire g17855;
wire II14948;
wire g18845;
wire II24409;
wire II37854;
wire II14808;
wire g24832;
wire II39071;
wire II31751;
wire g16527;
wire g28949;
wire II38101;
wire g12466;
wire g13999;
wire g4380;
wire II41123;
wire II37044;
wire g13117;
wire g9955;
wire g26682;
wire g5649;
wire g29262;
wire g24568;
wire g9113;
wire II27314;
wire g18999;
wire g4220;
wire g22340;
wire g22684;
wire II23153;
wire g8802;
wire g8523;
wire g28459;
wire g22100;
wire g28053;
wire g21522;
wire g13879;
wire g19471;
wire g22642;
wire g22383;
wire g26326;
wire g4951;
wire g8503;
wire g4456;
wire g25986;
wire II20431;
wire II20688;
wire g11784;
wire g25930;
wire g16880;
wire g16422;
wire g23244;
wire g23844;
wire g28287;
wire g10631;
wire g10182;
wire g29182;
wire II31586;
wire g10437;
wire g30440;
wire gbuf125;
wire g24421;
wire g30175;
wire II24036;
wire g4257;
wire II27755;
wire g16159;
wire g10724;
wire II36120;
wire g28373;
wire g30975;
wire g15332;
wire II24110;
wire g18886;
wire g13369;
wire g23081;
wire gbuf165;
wire g15245;
wire II17051;
wire II34707;
wire g29389;
wire II34764;
wire g9906;
wire II38644;
wire II21037;
wire g10010;
wire g18341;
wire g25445;
wire g5391;
wire g17091;
wire g24426;
wire II31814;
wire g13702;
wire g4749;
wire g13915;
wire g13320;
wire g28264;
wire g12039;
wire II21638;
wire g19124;
wire g29629;
wire g18432;
wire II30563;
wire II36162;
wire g16651;
wire g8945;
wire II30128;
wire II38831;
wire II14338;
wire II30092;
wire g30216;
wire g12079;
wire g22757;
wire g21420;
wire II21149;
wire g21425;
wire g26749;
wire II29040;
wire g30758;
wire g9441;
wire g23642;
wire g7354;
wire g5910;
wire g15259;
wire g9422;
wire II35539;
wire g5786;
wire g5807;
wire g18692;
wire g18899;
wire g24664;
wire II32067;
wire g29407;
wire g13601;
wire g13558;
wire g5233;
wire g26258;
wire g23229;
wire g28074;
wire g10059;
wire g28462;
wire g26960;
wire g30766;
wire g24240;
wire g28365;
wire g26257;
wire g25802;
wire II15986;
wire g17548;
wire g27522;
wire II24054;
wire g30723;
wire g11911;
wire g16182;
wire g13401;
wire II36052;
wire g18503;
wire g3522;
wire II24495;
wire II34296;
wire II18298;
wire g11701;
wire g28282;
wire g27976;
wire g30846;
wire g16938;
wire g26061;
wire g23222;
wire II21096;
wire g26307;
wire g26762;
wire II24679;
wire g21696;
wire g27140;
wire g13062;
wire g28310;
wire g9108;
wire g19711;
wire II35125;
wire g3710;
wire g27955;
wire II13804;
wire g21176;
wire g25163;
wire g24573;
wire II30221;
wire g8797;
wire g27354;
wire g23224;
wire g14936;
wire g20086;
wire II24639;
wire g18170;
wire II27338;
wire g26660;
wire g16831;
wire II34449;
wire g20346;
wire g24488;
wire g8576;
wire g17925;
wire II18734;
wire g5848;
wire II20398;
wire g13741;
wire g22164;
wire g26986;
wire g7815;
wire g4017;
wire II17009;
wire g28120;
wire g12291;
wire g19649;
wire g25208;
wire g27268;
wire g10281;
wire g8539;
wire g29437;
wire g10714;
wire g11872;
wire II34695;
wire g12895;
wire g8984;
wire g11656;
wire g22899;
wire g16673;
wire g12224;
wire g26082;
wire g28272;
wire g5836;
wire g23690;
wire g13174;
wire g20796;
wire g19261;
wire g4763;
wire II23943;
wire g19512;
wire gbuf49;
wire g24322;
wire g14685;
wire II18530;
wire g24314;
wire g10203;
wire II17681;
wire g17019;
wire g12352;
wire g27626;
wire g21163;
wire g15443;
wire g13343;
wire II31847;
wire g27324;
wire g6751;
wire g19160;
wire II19756;
wire g22384;
wire II39951;
wire g8918;
wire II34358;
wire II36465;
wire II30673;
wire g8396;
wire g25152;
wire g30749;
wire II34713;
wire g8031;
wire II19560;
wire g10430;
wire II31910;
wire g26429;
wire II38049;
wire II35404;
wire II14925;
wire II30735;
wire II32670;
wire g19299;
wire g18756;
wire II36609;
wire gbuf192;
wire g4561;
wire g20108;
wire II28524;
wire g21776;
wire g10011;
wire g15665;
wire g16906;
wire II26816;
wire g27746;
wire g12021;
wire II16700;
wire g12246;
wire g14885;
wire g28898;
wire g28420;
wire g27361;
wire g29794;
wire g17526;
wire g29221;
wire g28452;
wire g28335;
wire g16450;
wire g10393;
wire g21315;
wire g12100;
wire g20021;
wire gbuf66;
wire II19472;
wire g29320;
wire g26245;
wire g15604;
wire g9775;
wire g20525;
wire g22958;
wire g26675;
wire g20365;
wire g21243;
wire g5193;
wire g16575;
wire g17835;
wire g26186;
wire II37978;
wire g11691;
wire g27016;
wire g24128;
wire g20092;
wire g21086;
wire II20577;
wire g26581;
wire g18223;
wire g29259;
wire g10521;
wire g15808;
wire g4492;
wire II15922;
wire g21140;
wire g21730;
wire II24206;
wire g6014;
wire g19732;
wire II22752;
wire g27183;
wire II18674;
wire II36341;
wire II17854;
wire II37891;
wire g24589;
wire g13444;
wire II38139;
wire g29470;
wire II35106;
wire g23171;
wire g22988;
wire g29019;
wire II30230;
wire II35701;
wire II18578;
wire g19415;
wire g5129;
wire g30943;
wire II19961;
wire II25541;
wire g25996;
wire g22589;
wire g20752;
wire g29937;
wire g20816;
wire g15634;
wire II37047;
wire g21065;
wire g10250;
wire II22842;
wire II16811;
wire g18992;
wire g5148;
wire g7587;
wire g19315;
wire II39902;
wire g9585;
wire g26809;
wire g5280;
wire g27730;
wire g7855;
wire g17770;
wire g26300;
wire g5179;
wire g30327;
wire II32444;
wire II14104;
wire g10408;
wire g24224;
wire g8677;
wire II39369;
wire g26608;
wire II20421;
wire g24287;
wire g25146;
wire II13934;
wire g27905;
wire g13329;
wire g13399;
wire g27294;
wire g8427;
wire g25387;
wire II23584;
wire g12690;
wire g28677;
wire g5737;
wire g12121;
wire g17031;
wire g20473;
wire g30099;
wire II40203;
wire g5812;
wire g29243;
wire g14286;
wire g23778;
wire g24146;
wire g13867;
wire g19105;
wire g26959;
wire II40898;
wire g10494;
wire g25226;
wire g7534;
wire g7529;
wire g28400;
wire g3678;
wire g22191;
wire g11981;
wire g12125;
wire g22775;
wire g24068;
wire II36258;
wire g29346;
wire g20711;
wire g26571;
wire g17024;
wire g28187;
wire g5207;
wire II28994;
wire II26538;
wire g16803;
wire II17969;
wire g9367;
wire g26283;
wire g13360;
wire g24770;
wire II13655;
wire g12801;
wire g19869;
wire g5164;
wire II23475;
wire g17149;
wire II33188;
wire g25125;
wire g18650;
wire g29501;
wire g30284;
wire II40781;
wire g5050;
wire g10377;
wire g16082;
wire g22907;
wire g22876;
wire g26816;
wire II37358;
wire II39050;
wire g11538;
wire g11509;
wire g27783;
wire g5304;
wire g17738;
wire g30367;
wire g10214;
wire II34797;
wire g26618;
wire II32286;
wire II18214;
wire g8381;
wire g14280;
wire g16611;
wire g28919;
wire g30477;
wire g12931;
wire II32567;
wire II34077;
wire g17226;
wire g19054;
wire g28362;
wire g24331;
wire g18371;
wire II37822;
wire II26708;
wire g11160;
wire g9737;
wire II34080;
wire g20248;
wire g11994;
wire g4848;
wire g23782;
wire g12836;
wire g24207;
wire g29480;
wire g6974;
wire II25923;
wire g7664;
wire g28111;
wire g27482;
wire g28580;
wire g25752;
wire g28309;
wire g26012;
wire II39068;
wire II15532;
wire g21586;
wire II35049;
wire g24372;
wire g11330;
wire g25096;
wire g23550;
wire II18512;
wire g25288;
wire g20921;
wire g10238;
wire II30928;
wire g16985;
wire g14148;
wire II33580;
wire g26742;
wire g8937;
wire g11908;
wire g10295;
wire g4548;
wire II23083;
wire II37107;
wire g27566;
wire g27386;
wire g8756;
wire g13025;
wire g23857;
wire g30715;
wire g15385;
wire g21067;
wire g22283;
wire g21723;
wire g22461;
wire g10708;
wire g5656;
wire g24052;
wire g29574;
wire II38872;
wire g22319;
wire II15806;
wire g13195;
wire g8000;
wire g27997;
wire II15850;
wire g21558;
wire g30104;
wire g24582;
wire g21822;
wire g3806;
wire g28704;
wire II23143;
wire g11795;
wire II38250;
wire g28044;
wire g21467;
wire g7338;
wire g15553;
wire g23551;
wire g26737;
wire g20928;
wire II25856;
wire g21107;
wire II34946;
wire g16016;
wire II14763;
wire II39631;
wire g5551;
wire g27297;
wire g22694;
wire g15262;
wire g23277;
wire g19209;
wire g12430;
wire g24523;
wire g21871;
wire g14183;
wire g17718;
wire g25412;
wire g29112;
wire g14795;
wire g5939;
wire II13896;
wire g4552;
wire g26157;
wire gbuf187;
wire g23872;
wire g29300;
wire g24341;
wire II36960;
wire g26645;
wire g25588;
wire g26508;
wire II22524;
wire g24754;
wire II32547;
wire g5057;
wire g7879;
wire g8517;
wire g30308;
wire g26719;
wire g29686;
wire g29097;
wire g26498;
wire g22887;
wire g24880;
wire II29351;
wire g20447;
wire g23359;
wire II26667;
wire g20971;
wire II32871;
wire g23557;
wire II39638;
wire g20570;
wire g20241;
wire II30284;
wire g14431;
wire g30504;
wire g30072;
wire II37804;
wire g6519;
wire g19902;
wire g6100;
wire II21364;
wire g23588;
wire II28155;
wire g25378;
wire II27391;
wire g10329;
wire g21118;
wire g24432;
wire g21123;
wire II34505;
wire g11865;
wire g26657;
wire g19941;
wire g5622;
wire g17051;
wire II15651;
wire g19796;
wire g18369;
wire II28162;
wire g21878;
wire g22247;
wire II28174;
wire II26396;
wire II23712;
wire g5775;
wire g24405;
wire g24656;
wire g16507;
wire g14641;
wire g11271;
wire II14618;
wire II34124;
wire g28863;
wire II36426;
wire II14605;
wire II17774;
wire g29395;
wire g27548;
wire g24904;
wire II39800;
wire II40128;
wire g23953;
wire g13166;
wire g21455;
wire g11410;
wire g25233;
wire g7712;
wire g29142;
wire g4211;
wire g22080;
wire II30725;
wire g25013;
wire II29375;
wire II18452;
wire II37295;
wire g28163;
wire g11737;
wire g8931;
wire g26730;
wire II22918;
wire II15543;
wire g12370;
wire g10678;
wire g15877;
wire g25859;
wire g29361;
wire II38474;
wire g18796;
wire g26635;
wire g29755;
wire II14577;
wire g29609;
wire II38496;
wire g28174;
wire g16264;
wire g25400;
wire II27822;
wire g29317;
wire II16015;
wire II32961;
wire II31499;
wire g26613;
wire II19208;
wire II26357;
wire g30285;
wire g5953;
wire II34983;
wire g27033;
wire g27023;
wire II29310;
wire II40618;
wire g13184;
wire g27707;
wire II25809;
wire g14028;
wire g28223;
wire g24443;
wire g10510;
wire II18277;
wire g21932;
wire g24412;
wire g5604;
wire g17255;
wire g27962;
wire g13463;
wire g23860;
wire g23160;
wire II26676;
wire g20116;
wire II38352;
wire g30293;
wire g20085;
wire g16483;
wire g19190;
wire II32988;
wire g5895;
wire g25732;
wire g25513;
wire g24472;
wire II39089;
wire g15094;
wire g17151;
wire g22999;
wire g12504;
wire II26500;
wire II37912;
wire II27203;
wire g17882;
wire g27814;
wire g18414;
wire g13499;
wire g29281;
wire g28567;
wire g13218;
wire g28340;
wire g23900;
wire g27759;
wire g25052;
wire g5408;
wire g11880;
wire II38483;
wire g11007;
wire g8564;
wire g16107;
wire II26545;
wire g24558;
wire g19787;
wire g10650;
wire II22763;
wire g22139;
wire g19970;
wire II23217;
wire gbuf210;
wire II30829;
wire II28485;
wire II33526;
wire gbuf83;
wire g29303;
wire g4427;
wire II19557;
wire g26396;
wire g19842;
wire g24004;
wire II36867;
wire g30647;
wire g13421;
wire II17945;
wire g19204;
wire II13913;
wire II36141;
wire g10044;
wire II35923;
wire g5662;
wire II35476;
wire g5389;
wire g12851;
wire g24604;
wire II29408;
wire g30131;
wire g25530;
wire g16702;
wire g24551;
wire g23233;
wire II34063;
wire g29881;
wire II19488;
wire g29555;
wire II23208;
wire g12008;
wire g30728;
wire g29398;
wire g24280;
wire g28416;
wire g25139;
wire II37920;
wire g16187;
wire g6212;
wire g21414;
wire g5951;
wire g12142;
wire g9112;
wire g9306;
wire g4507;
wire II22683;
wire II33801;
wire g25073;
wire II18108;
wire g30263;
wire g21023;
wire g9419;
wire g8654;
wire g13095;
wire g10166;
wire g5746;
wire II23345;
wire g23771;
wire g13427;
wire g18720;
wire g29974;
wire II30185;
wire II38999;
wire g23910;
wire g27775;
wire II38716;
wire II21497;
wire II20604;
wire g27413;
wire g28681;
wire g25443;
wire g26168;
wire g3237;
wire g16014;
wire g12429;
wire g19026;
wire g9123;
wire II29690;
wire II37330;
wire g19722;
wire gbuf24;
wire g26295;
wire g26407;
wire g11382;
wire g10617;
wire g8665;
wire g29663;
wire g10548;
wire g5504;
wire g4725;
wire g23726;
wire g25426;
wire g5627;
wire g24704;
wire g24254;
wire g18655;
wire g25776;
wire g20388;
wire g15127;
wire g26386;
wire II16544;
wire g23432;
wire g7766;
wire II13152;
wire g15353;
wire g10107;
wire II27491;
wire g26144;
wire g8502;
wire g12955;
wire g23531;
wire g18810;
wire II21523;
wire g23158;
wire II25092;
wire g22177;
wire g10331;
wire g13418;
wire II22702;
wire II26320;
wire g11763;
wire g17433;
wire g19227;
wire II19321;
wire g10112;
wire II23863;
wire II33374;
wire g10866;
wire II36936;
wire g24530;
wire II36367;
wire g4282;
wire II21936;
wire g30336;
wire g19288;
wire II23588;
wire II33825;
wire g30773;
wire g9807;
wire g26415;
wire g20341;
wire g19747;
wire II27426;
wire g16324;
wire g28983;
wire g21598;
wire II29212;
wire II26134;
wire g7460;
wire II14599;
wire g5819;
wire g26798;
wire g24512;
wire g29764;
wire II24923;
wire g17796;
wire g9080;
wire g8059;
wire II27002;
wire II21446;
wire g24111;
wire II16469;
wire II36696;
wire g5098;
wire II25554;
wire II29566;
wire II15481;
wire g18539;
wire g26221;
wire g8255;
wire g30011;
wire g10968;
wire g13147;
wire g11947;
wire II38258;
wire II23670;
wire g19444;
wire g27330;
wire g23211;
wire II33219;
wire g19593;
wire g26756;
wire g28292;
wire g26690;
wire g18894;
wire g13492;
wire g6777;
wire g16062;
wire II23027;
wire g29511;
wire g15700;
wire II18085;
wire g19352;
wire g8587;
wire g17182;
wire g14321;
wire g23562;
wire g20103;
wire II37125;
wire g12650;
wire g13901;
wire II25872;
wire g25947;
wire g25099;
wire II32295;
wire g18957;
wire g12421;
wire g15429;
wire g18914;
wire g11327;
wire g26701;
wire g28732;
wire g22699;
wire II19552;
wire g30964;
wire g15458;
wire g22590;
wire g20336;
wire II31739;
wire g28206;
wire g27337;
wire g7475;
wire g15561;
wire g15888;
wire g19131;
wire II32439;
wire g28357;
wire g26030;
wire g28488;
wire g10226;
wire g18929;
wire II27240;
wire g28707;
wire g26935;
wire II18166;
wire II18157;
wire II30991;
wire g4324;
wire g21521;
wire g28747;
wire g8912;
wire g9056;
wire g24466;
wire g30314;
wire g13103;
wire II39773;
wire g29692;
wire II27131;
wire g23207;
wire g29416;
wire g10644;
wire II29001;
wire g18634;
wire g27743;
wire g23603;
wire II17727;
wire g12268;
wire g19533;
wire II24437;
wire II38018;
wire II38713;
wire gbuf96;
wire g22664;
wire g21376;
wire II39534;
wire g4929;
wire g20137;
wire II37161;
wire g19880;
wire g24303;
wire g11935;
wire g16813;
wire g13528;
wire g24461;
wire g22936;
wire g9096;
wire g16212;
wire g25160;
wire g13072;
wire g7614;
wire g16283;
wire g27122;
wire g26638;
wire gbuf12;
wire II14535;
wire g13292;
wire g22005;
wire g5110;
wire II35355;
wire II23817;
wire g29523;
wire g15439;
wire g24408;
wire g9076;
wire gbuf197;
wire II20523;
wire g12059;
wire g17117;
wire II30137;
wire g9464;
wire g23743;
wire g29411;
wire II24894;
wire g24103;
wire g22700;
wire II14888;
wire g10986;
wire g25793;
wire II18197;
wire g13892;
wire g19540;
wire g9391;
wire g5593;
wire g27761;
wire II19342;
wire g26672;
wire II23845;
wire II28152;
wire g6305;
wire g29751;
wire g26067;
wire g17436;
wire g30802;
wire g4104;
wire g5736;
wire g22724;
wire g22397;
wire II16221;
wire II30107;
wire g23146;
wire g30614;
wire g26586;
wire g10351;
wire g30863;
wire II35153;
wire g10817;
wire g21954;
wire g9607;
wire g16043;
wire g24370;
wire g19212;
wire II21580;
wire g10076;
wire g21309;
wire g5341;
wire g4683;
wire g19930;
wire g24591;
wire II26476;
wire g16385;
wire g4147;
wire g18865;
wire g23765;
wire g22608;
wire g8009;
wire g23923;
wire g7721;
wire II18629;
wire g22519;
wire g15197;
wire g27161;
wire g16442;
wire g28449;
wire g24882;
wire g14613;
wire g19811;
wire g28157;
wire II36563;
wire g30912;
wire g21886;
wire II33361;
wire g5858;
wire g18036;
wire g21735;
wire II25692;
wire g15221;
wire g23100;
wire g23591;
wire g30686;
wire g11490;
wire g12907;
wire g13348;
wire II36246;
wire g11777;
wire II16252;
wire g10629;
wire g15115;
wire g9857;
wire g4994;
wire g23308;
wire g19418;
wire g30979;
wire II38154;
wire g23891;
wire II37386;
wire g19383;
wire II37650;
wire g30786;
wire g22647;
wire g23730;
wire g27166;
wire g21041;
wire II25742;
wire g24687;
wire II18217;
wire g18903;
wire II13366;
wire g20007;
wire g26820;
wire g24675;
wire g1942;
wire g27854;
wire II21531;
wire II26985;
wire g20598;
wire g29536;
wire g30115;
wire g5762;
wire g18668;
wire II22557;
wire g14570;
wire II36714;
wire II17156;
wire g30373;
wire II18560;
wire II36653;
wire g8808;
wire g24211;
wire g10800;
wire g5873;
wire g10921;
wire g21093;
wire g25241;
wire g24115;
wire g25870;
wire g9132;
wire II30757;
wire g8824;
wire g25085;
wire II18491;
wire g25981;
wire II18229;
wire II28521;
wire g4254;
wire g11966;
wire g13787;
wire II36354;
wire g23660;
wire g15922;
wire II27077;
wire II21998;
wire g20577;
wire II17734;
wire II25456;
wire g28713;
wire II37514;
wire g7718;
wire g9965;
wire g16996;
wire g20219;
wire II40119;
wire g10659;
wire g28006;
wire g14959;
wire g17357;
wire g13646;
wire II13910;
wire g9958;
wire g18278;
wire g29185;
wire II32511;
wire g23720;
wire g16010;
wire g24548;
wire g8475;
wire g22376;
wire II31031;
wire g17627;
wire II13901;
wire g16251;
wire g14027;
wire g12493;
wire g17394;
wire II24494;
wire g19786;
wire g29263;
wire II15577;
wire g11624;
wire g4532;
wire g7833;
wire g29608;
wire g26597;
wire g13041;
wire g11690;
wire g29368;
wire g17741;
wire g23381;
wire g19890;
wire g13299;
wire g26954;
wire g8242;
wire g28271;
wire g20621;
wire g13300;
wire g17449;
wire g5044;
wire II28754;
wire II24753;
wire g23388;
wire g15836;
wire II13182;
wire g28214;
wire g4085;
wire g20561;
wire g14471;
wire g6438;
wire II30878;
wire II20458;
wire g8579;
wire II25612;
wire g28442;
wire g13010;
wire II37868;
wire II31162;
wire g21921;
wire g20268;
wire g23200;
wire II40429;
wire g30879;
wire g17234;
wire g4857;
wire g23682;
wire II29203;
wire g23427;
wire g12052;
wire II38594;
wire II15493;
wire g24468;
wire g10479;
wire g16935;
wire g7420;
wire g19515;
wire g12152;
wire II34230;
wire g27054;
wire II23076;
wire g13675;
wire II24545;
wire g19016;
wire g23180;
wire g30857;
wire II31451;
wire II23893;
wire g29914;
wire II18632;
wire g24736;
wire g11373;
wire II18611;
wire g28892;
wire g11866;
wire g17383;
wire g30021;
wire g16778;
wire g29727;
wire II15918;
wire g30841;
wire g29274;
wire g24874;
wire g7583;
wire g21169;
wire g13370;
wire g18490;
wire g22343;
wire g20842;
wire II32164;
wire g10809;
wire II40730;
wire II36536;
wire II25044;
wire g26988;
wire II17030;
wire gbuf175;
wire II24078;
wire g24455;
wire g29154;
wire II23046;
wire g25047;
wire g22776;
wire g26214;
wire II29918;
wire g17950;
wire II29963;
wire II28503;
wire g18960;
wire g22745;
wire g30081;
wire II21897;
wire g25362;
wire g26778;
wire II13218;
wire g13677;
wire g9781;
wire g17541;
wire g27264;
wire g23713;
wire g16233;
wire g10711;
wire II18013;
wire g8785;
wire II14550;
wire II22912;
wire g12914;
wire II21992;
wire g20058;
wire g28385;
wire g16964;
wire g12221;
wire g5878;
wire II37092;
wire g12997;
wire g30002;
wire g12326;
wire II38453;
wire g18875;
wire g4570;
wire g20049;
wire g23030;
wire g28107;
wire II20634;
wire g3981;
wire g29111;
wire II36741;
wire g30807;
wire g25217;
wire g12814;
wire g11255;
wire II31625;
wire II20863;
wire II25800;
wire g22107;
wire g24843;
wire g10302;
wire g8760;
wire g30353;
wire II37584;
wire g20877;
wire g5929;
wire g5759;
wire g21667;
wire g5740;
wire II40775;
wire g15812;
wire g12091;
wire g20315;
wire g8417;
wire g25348;
wire g8688;
wire g27129;
wire g22306;
wire g30277;
wire g28239;
wire g15338;
wire g19062;
wire g13622;
wire II35886;
wire II27972;
wire g25877;
wire g27234;
wire g30572;
wire II39038;
wire g5095;
wire g23314;
wire II39997;
wire g16313;
wire II36253;
wire g24925;
wire g14606;
wire II23625;
wire g10291;
wire g18623;
wire g27671;
wire g11588;
wire g13880;
wire g10821;
wire g11210;
wire II40751;
wire g20323;
wire g17192;
wire g23190;
wire g29191;
wire II32357;
wire g10288;
wire g17059;
wire g10689;
wire g12477;
wire g20062;
wire g27493;
wire g29236;
wire g6636;
wire g19172;
wire g14565;
wire II23513;
wire g20015;
wire g25109;
wire II31859;
wire II30113;
wire g17229;
wire II38515;
wire g17097;
wire g25187;
wire g12939;
wire II20703;
wire g24347;
wire II40313;
wire g10663;
wire g11794;
wire g12069;
wire g29139;
wire g18946;
wire g22736;
wire g23892;
wire g29788;
wire g4573;
wire g14249;
wire gbuf7;
wire g25314;
wire g26689;
wire II17061;
wire g18953;
wire g15783;
wire g30517;
wire g13156;
wire g13378;
wire g16866;
wire II29990;
wire II21796;
wire g22661;
wire g20977;
wire II20359;
wire g16468;
wire g9822;
wire II28357;
wire II35834;
wire II34388;
wire g5697;
wire g11678;
wire II26285;
wire g11392;
wire g18833;
wire g10928;
wire g11929;
wire g20557;
wire g29425;
wire II25423;
wire g19278;
wire g27631;
wire g24888;
wire g4107;
wire g11277;
wire II20652;
wire g13200;
wire II25644;
wire g8378;
wire g21988;
wire g29491;
wire g22210;
wire g4118;
wire g13079;
wire g13322;
wire II20813;
wire g30643;
wire g26887;
wire g7891;
wire II31685;
wire g30129;
wire g20437;
wire g25333;
wire g8071;
wire g14171;
wire g18920;
wire g21651;
wire II18653;
wire II13928;
wire II14654;
wire g25488;
wire g8842;
wire g19159;
wire g7806;
wire II35708;
wire g29455;
wire II37632;
wire g27045;
wire II23445;
wire g24819;
wire g26004;
wire g23084;
wire g5922;
wire g21001;
wire gbuf41;
wire g20717;
wire g17001;
wire g8990;
wire g25369;
wire II17125;
wire g20146;
wire II40883;
wire II29653;
wire g24957;
wire II31124;
wire II33479;
wire g23792;
wire g26106;
wire g23199;
wire g25886;
wire g20605;
wire g23344;
wire II26198;
wire g27325;
wire g6205;
wire g27541;
wire g25145;
wire g27513;
wire g8215;
wire g18763;
wire II40661;
wire II25334;
wire g9506;
wire g16300;
wire g19271;
wire g24800;
wire II17106;
wire g18836;
wire g18598;
wire g15793;
wire g11919;
wire g27098;
wire II24725;
wire g17399;
wire g11503;
wire g29457;
wire g19852;
wire g30225;
wire g23189;
wire g19594;
wire g26530;
wire gbuf19;
wire g17825;
wire g7195;
wire g8317;
wire II21868;
wire g12062;
wire g28690;
wire g29545;
wire II28235;
wire g19256;
wire II14502;
wire II40086;
wire g25008;
wire g28785;
wire g22208;
wire g10449;
wire g29064;
wire g28814;
wire II35512;
wire II24399;
wire g17959;
wire g21403;
wire g5659;
wire g27551;
wire II24196;
wire g20061;
wire g21788;
wire II15677;
wire g6232;
wire g26981;
wire g22215;
wire gbuf54;
wire g29128;
wire g26625;
wire g10442;
wire g16254;
wire II31556;
wire g14497;
wire g15453;
wire g26458;
wire g30587;
wire g18297;
wire g28788;
wire II33352;
wire g4578;
wire II14343;
wire g28609;
wire g5852;
wire g16239;
wire g25972;
wire g19106;
wire II24187;
wire g29953;
wire g24416;
wire g20399;
wire g30108;
wire II18641;
wire g11581;
wire g28016;
wire g8076;
wire g13755;
wire g11510;
wire g21808;
wire II25561;
wire gbuf206;
wire g19950;
wire g30923;
wire g9887;
wire g10589;
wire g19147;
wire g23482;
wire g28883;
wire g30040;
wire g28323;
wire g19701;
wire g15822;
wire II33810;
wire g8543;
wire II24340;
wire g27144;
wire g21198;
wire g28726;
wire g25386;
wire g20283;
wire g16459;
wire g18302;
wire II30320;
wire g23573;
wire II13980;
wire II32460;
wire g21855;
wire g27384;
wire g13502;
wire g29985;
wire g14290;
wire g3996;
wire g18881;
wire II40578;
wire g7706;
wire g28733;
wire g29446;
wire g29254;
wire g17172;
wire g10500;
wire g7730;
wire g22234;
wire g4879;
wire II31691;
wire g29569;
wire gbuf162;
wire g23637;
wire g6081;
wire g19357;
wire g29441;
wire g13536;
wire g20303;
wire II24640;
wire II15565;
wire II36479;
wire g5866;
wire II16027;
wire g4655;
wire g20374;
wire g23017;
wire II29948;
wire g27036;
wire II13161;
wire g27240;
wire II20517;
wire g27938;
wire II24318;
wire g19719;
wire g29869;
wire g10156;
wire g27197;
wire g20624;
wire g12433;
wire g9746;
wire II28115;
wire II38450;
wire g26090;
wire g21517;
wire II17043;
wire g8748;
wire g8177;
wire II29712;
wire II37986;
wire g22259;
wire g11803;
wire g9371;
wire g10354;
wire g5700;
wire g18604;
wire g21654;
wire g28458;
wire g23266;
wire g22530;
wire g21514;
wire g13635;
wire g27572;
wire g5830;
wire II18761;
wire II22651;
wire g15829;
wire g5081;
wire g24440;
wire g16712;
wire g22563;
wire g27079;
wire g19565;
wire g11932;
wire g20089;
wire g20288;
wire II32193;
wire g4504;
wire g15994;
wire g8194;
wire g26031;
wire g9939;
wire II35446;
wire g11799;
wire g9006;
wire g10065;
wire II18584;
wire g15950;
wire g29947;
wire g8627;
wire g24498;
wire g16336;
wire II15946;
wire II36876;
wire II39243;
wire g24095;
wire g20330;
wire g28967;
wire g25327;
wire g10458;
wire g30885;
wire II29049;
wire g24175;
wire II20694;
wire g10534;
wire g21329;
wire g21380;
wire g3337;
wire g24271;
wire g14609;
wire g21494;
wire g22428;
wire II30614;
wire II39818;
wire g13000;
wire g23944;
wire II17370;
wire II21723;
wire g25192;
wire g24380;
wire g21011;
wire g18314;
wire II27257;
wire g20080;
wire g27942;
wire g28097;
wire II18103;
wire II34650;
wire g15699;
wire g5072;
wire II23836;
wire g20486;
wire g22054;
wire g27594;
wire II32402;
wire g23286;
wire g22163;
wire g15803;
wire g11825;
wire II30797;
wire g25156;
wire g12212;
wire II32597;
wire II28726;
wire g24327;
wire g24470;
wire g19035;
wire g17446;
wire g30894;
wire g16907;
wire g19171;
wire g5382;
wire g30951;
wire g26692;
wire g14773;
wire g24114;
wire g20456;
wire II32669;
wire g14039;
wire g18986;
wire g28306;
wire II17685;
wire g5887;
wire g21396;
wire g29420;
wire g25320;
wire II37059;
wire g17471;
wire II16065;
wire g12972;
wire II18542;
wire g8569;
wire g11264;
wire g21158;
wire g23285;
wire II29603;
wire g27988;
wire g4079;
wire g23617;
wire g24278;
wire II26966;
wire g6039;
wire II38321;
wire g11638;
wire II35883;
wire g9064;
wire g12537;
wire g29331;
wire II14973;
wire g21594;
wire g26793;
wire g14252;
wire g29993;
wire g10612;
wire II33246;
wire g20538;
wire g21627;
wire II20493;
wire g16595;
wire g27027;
wire g11742;
wire g11098;
wire II35036;
wire II39339;
wire g23827;
wire II14857;
wire g16113;
wire II13953;
wire g24479;
wire g29758;
wire g22790;
wire II28061;
wire g13110;
wire II18265;
wire g27020;
wire g30952;
wire II38626;
wire g3941;
wire II32889;
wire g27969;
wire g26605;
wire II18241;
wire g22728;
wire g29657;
wire g20442;
wire g22490;
wire g22881;
wire g26261;
wire II21933;
wire II32140;
wire g12859;
wire II27083;
wire g13922;
wire II39916;
wire II21274;
wire g25515;
wire g13856;
wire g17563;
wire g16003;
wire g17530;
wire g26548;
wire g8203;
wire g28250;
wire g22620;
wire g30774;
wire II34032;
wire g29775;
wire g4082;
wire g25177;
wire g9116;
wire II19507;
wire g7541;
wire g29373;
wire g19468;
wire II20032;
wire g23630;
wire g18619;
wire g26291;
wire g21687;
wire g6675;
wire g27249;
wire g5508;
wire g26471;
wire g27225;
wire g23291;
wire g19450;
wire g26906;
wire g16344;
wire g24809;
wire II19500;
wire g22556;
wire g3247;
wire g25141;
wire g23087;
wire g13394;
wire g11179;
wire g23230;
wire g9819;
wire II25783;
wire g15859;
wire g8484;
wire gbuf215;
wire g29770;
wire II18025;
wire g13207;
wire II14424;
wire g10431;
wire g20397;
wire II23878;
wire g25281;
wire g10541;
wire g12251;
wire g12498;
wire g27912;
wire II17709;
wire gbuf39;
wire g13247;
wire g17579;
wire g12825;
wire II29456;
wire g15739;
wire II37277;
wire g26789;
wire g14024;
wire II23992;
wire II31253;
wire g27716;
wire II26348;
wire g4351;
wire g18866;
wire g24143;
wire g29808;
wire g28838;
wire g24389;
wire II22542;
wire g20898;
wire g21196;
wire g8512;
wire g7691;
wire II40149;
wire g23461;
wire II27140;
wire II25763;
wire g30465;
wire II35376;
wire g28046;
wire g11592;
wire g30276;
wire g4315;
wire g9816;
wire II38881;
wire g23544;
wire II26934;
wire g27959;
wire g23360;
wire II29183;
wire II34029;
wire g24789;
wire g18011;
wire g17275;
wire g30785;
wire g30818;
wire g26724;
wire g4734;
wire g16023;
wire II39340;
wire g18395;
wire II31088;
wire g5663;
wire g12445;
wire g29147;
wire g21143;
wire g26516;
wire g28433;
wire g10875;
wire g13327;
wire g22361;
wire g29849;
wire II13925;
wire g27496;
wire g29547;
wire g25711;
wire II23430;
wire II39414;
wire g24768;
wire g24526;
wire II24006;
wire II34997;
wire g15109;
wire II36296;
wire g29381;
wire II38003;
wire g19752;
wire II27170;
wire II27308;
wire II16092;
wire g18842;
wire g21260;
wire II20574;
wire g26972;
wire g19553;
wire g23721;
wire g26315;
wire g27682;
wire II38181;
wire g27102;
wire g17422;
wire II29872;
wire g8015;
wire g10691;
wire II29246;
wire g19772;
wire g23125;
wire g11997;
wire g23508;
wire g8433;
wire g24865;
wire g25203;
wire g4275;
wire II30766;
wire g21138;
wire gbuf113;
wire g18794;
wire II37110;
wire g6018;
wire g20951;
wire g22335;
wire g13614;
wire g10898;
wire g24501;
wire g25026;
wire g10973;
wire g23766;
wire g13788;
wire g8949;
wire II37119;
wire g6139;
wire g11728;
wire g21290;
wire g29170;
wire g5415;
wire g19523;
wire g20298;
wire g26404;
wire II32308;
wire II17884;
wire II40542;
wire g28772;
wire g21120;
wire g23149;
wire g27307;
wire gbuf158;
wire g18639;
wire g21470;
wire II40521;
wire g24508;
wire g9641;
wire g13436;
wire g30811;
wire II32626;
wire g12114;
wire g13547;
wire g5399;
wire g9128;
wire g5771;
wire g26568;
wire g28986;
wire II25123;
wire g21078;
wire g24751;
wire g19308;
wire g8483;
wire g15660;
wire g23420;
wire g18351;
wire g27721;
wire g4159;
wire II37939;
wire II40555;
wire g26160;
wire g19057;
wire g15254;
wire II32137;
wire g22060;
wire II39386;
wire g24437;
wire g5298;
wire II19598;
wire g27805;
wire g28347;
wire g17049;
wire II35750;
wire g29217;
wire g25560;
wire II34020;
wire g15317;
wire g16128;
wire g23777;
wire g15899;
wire g22803;
wire g3954;
wire g22844;
wire II20407;
wire g15234;
wire g28928;
wire g7575;
wire g10314;
wire II40913;
wire g19680;
wire g28411;
wire g30054;
wire II40242;
wire g22784;
wire g21962;
wire g20629;
wire g30487;
wire g9099;
wire g5940;
wire II36126;
wire g26864;
wire II30182;
wire g23401;
wire g19871;
wire g21816;
wire g9812;
wire g30837;
wire g24560;
wire g22189;
wire g8513;
wire g16025;
wire g11542;
wire gbuf104;
wire II16462;
wire g28217;
wire g11838;
wire g8561;
wire g3722;
wire g22311;
wire g25306;
wire g8693;
wire g10744;
wire II35076;
wire g25236;
wire g23581;
wire g4894;
wire g22711;
wire g27451;
wire g27151;
wire g11974;
wire g17314;
wire II31874;
wire g22506;
wire g10664;
wire g18781;
wire II25162;
wire II23348;
wire g29197;
wire g24334;
wire g21862;
wire g26810;
wire g27203;
wire g24391;
wire g26233;
wire g26017;
wire g8851;
wire II36362;
wire g17735;
wire g15904;
wire g5278;
wire g14186;
wire II33205;
wire II32860;
wire g9662;
wire II40260;
wire g30323;
wire g20982;
wire g25903;
wire II24438;
wire g27727;
wire g5366;
wire II30371;
wire g28649;
wire g15850;
wire II15839;
wire g21949;
wire g28021;
wire II30065;
wire g29803;
wire g15519;
wire g17341;
wire g28114;
wire g29933;
wire g8867;
wire g21103;
wire II33145;
wire g30349;
wire II33554;
wire g14118;
wire II28047;
wire g10671;
wire g30391;
wire g29688;
wire g24364;
wire g12084;
wire g19911;
wire II30344;
wire g28653;
wire g29560;
wire g7862;
wire g11735;
wire g6024;
wire II19747;
wire g30536;
wire g14831;
wire g26995;
wire g21363;
wire g4175;
wire II40215;
wire g27343;
wire g27373;
wire g15047;
wire g21572;
wire II39377;
wire g10434;
wire g30562;
wire g14725;
wire g5614;
wire g9968;
wire II18962;
wire g16463;
wire g8900;
wire g21344;
wire g5611;
wire II18563;
wire II29274;
wire II28479;
wire g5334;
wire g23303;
wire g22359;
wire g18647;
wire g16222;
wire II29797;
wire g5634;
wire II14621;
wire g8527;
wire g26334;
wire g19854;
wire g25685;
wire g4870;
wire g30335;
wire g7649;
wire g24890;
wire II21289;
wire II27062;
wire g24939;
wire g11493;
wire g20833;
wire g26801;
wire g19239;
wire II24576;
wire g18109;
wire g8101;
wire g5156;
wire g4888;
wire g30496;
wire g21320;
wire g26622;
wire II19722;
wire II25280;
wire II14442;
wire g8328;
wire g30705;
wire g12373;
wire g24294;
wire g12646;
wire g11526;
wire g28179;
wire g11036;
wire II29509;
wire II23132;
wire g20217;
wire g5631;
wire g11578;
wire II26923;
wire II30938;
wire II16993;
wire g29356;
wire II16457;
wire II14734;
wire g13565;
wire II29223;
wire g8829;
wire g15064;
wire g25129;
wire g28475;
wire g5315;
wire g28867;
wire g25579;
wire II38275;
wire II27684;
wire g29202;
wire g27088;
wire g25449;
wire II30875;
wire g23848;
wire g13706;
wire g10514;
wire II13931;
wire II34683;
wire g25934;
wire II23209;
wire g29625;
wire g23643;
wire II26599;
wire II25165;
wire g27131;
wire g4483;
wire g29406;
wire g11571;
wire g27917;
wire II28159;
wire g30781;
wire II30917;
wire g11941;
wire g11915;
wire II21398;
wire g27984;
wire g9779;
wire II28107;
wire g30753;
wire g26529;
wire g23093;
wire g8181;
wire g29223;
wire g4591;
wire g26766;
wire g11780;
wire II23034;
wire g16539;
wire g19933;
wire g29637;
wire g9890;
wire g5803;
wire g29500;
wire II30623;
wire g29086;
wire II34782;
wire II31565;
wire g3240;
wire g25205;
wire II34425;
wire g8312;
wire g28465;
wire II27318;
wire g11607;
wire g13183;
wire g30453;
wire g26026;
wire g23492;
wire g27622;
wire g23888;
wire g23225;
wire g13058;
wire II21747;
wire II21426;
wire II40236;
wire II26819;
wire II24278;
wire g22690;
wire II24158;
wire g15652;
wire II23472;
wire II23084;
wire II38704;
wire g28644;
wire II22945;
wire g9117;
wire g13263;
wire g16570;
wire g10838;
wire g30868;
wire g15393;
wire g17294;
wire g19266;
wire g26664;
wire g4806;
wire g19627;
wire g12781;
wire g27006;
wire g30529;
wire g9104;
wire g28668;
wire II14516;
wire g3617;
wire g29798;
wire g7391;
wire g14000;
wire g27864;
wire g23008;
wire gbuf122;
wire g8594;
wire II37572;
wire g27136;
wire g22681;
wire g22129;
wire g13196;
wire g7845;
wire II31727;
wire g28893;
wire g4026;
wire gbuf129;
wire g19298;
wire g15682;
wire g25850;
wire II18599;
wire g28286;
wire g5426;
wire g26964;
wire g29747;
wire g20418;
wire g13998;
wire g20367;
wire g5769;
wire g30638;
wire g13405;
wire g18626;
wire g25111;
wire g19975;
wire g29505;
wire g4452;
wire g17859;
wire g3304;
wire g26226;
wire g19983;
wire g8572;
wire g25890;
wire g5204;
wire II32325;
wire g7085;
wire g4829;
wire g30138;
wire II34986;
wire II31071;
wire g30406;
wire g26842;
wire II16987;
wire II13116;
wire g16007;
wire g16349;
wire g11859;
wire g20498;
wire g30171;
wire g26897;
wire g4032;
wire g19826;
wire g24422;
wire II18784;
wire II30257;
wire II38486;
wire g29385;
wire g22403;
wire g28958;
wire II17159;
wire II22755;
wire II35844;
wire g7923;
wire g5021;
wire II30038;
wire g17688;
wire g25016;
wire g25779;
wire g11988;
wire II38746;
wire II26871;
wire II17209;
wire g9921;
wire g21760;
wire g15804;
wire g19296;
wire g29134;
wire II25840;
wire g11054;
wire g21421;
wire g22914;
wire g12249;
wire g18617;
wire g13364;
wire g17442;
wire g25258;
wire g10517;
wire g5904;
wire II15484;
wire g16291;
wire g12899;
wire g30690;
wire II19289;
wire g28630;
wire II20462;
wire II37005;
wire g13088;
wire II36656;
wire g24708;
wire g24299;
wire g12025;
wire g22026;
wire g25989;
wire II40571;
wire g29324;
wire g22380;
wire g4357;
wire g24028;
wire g29651;
wire g13510;
wire II37481;
wire II19826;
wire g30918;
wire g23329;
wire g20647;
wire g19258;
wire g22543;
wire II31820;
wire g28194;
wire g13440;
wire g23575;
wire II36618;
wire II35551;
wire g30874;
wire g25703;
wire g25569;
wire g30911;
wire g12035;
wire g26649;
wire g21359;
wire g22668;
wire II18551;
wire g28124;
wire II21841;
wire g26555;
wire g24081;
wire II14590;
wire g5833;
wire II20682;
wire g27992;
wire II32133;
wire g19783;
wire g28247;
wire g9745;
wire g26086;
wire g23025;
wire g19640;
wire g7819;
wire II32198;
wire g27588;
wire g23830;
wire g19689;
wire g16162;
wire g29650;
wire g29971;
wire g30906;
wire II26535;
wire g30566;
wire g27951;
wire g13178;
wire g30247;
wire g25992;
wire g27910;
wire II23983;
wire g4626;
wire II37662;
wire II14637;
wire II20049;
wire II16942;
wire g20242;
wire g24585;
wire g19322;
wire g25962;
wire g23858;
wire g8286;
wire II23733;
wire g11398;
wire g5190;
wire g13479;
wire g22537;
wire II21688;
wire g28637;
wire g12228;
wire g25056;
wire g27273;
wire g25700;
wire II25210;
wire g26746;
wire g8459;
wire g10486;
wire II30101;
wire g22069;
wire II40982;
wire g19319;
wire g4016;
wire g25483;
wire g11123;
wire g30095;
wire g24326;
wire g24258;
wire g18590;
wire II27293;
wire II32478;
wire g20505;
wire II29503;
wire g6020;
wire g26187;
wire g23864;
wire g6047;
wire gbuf21;
wire g28276;
wire g17774;
wire g20423;
wire II17881;
wire g29403;
wire g26424;
wire g5411;
wire g29768;
wire g30551;
wire g22093;
wire g11011;
wire II24285;
wire g17520;
wire g22984;
wire g28424;
wire g24290;
wire II29981;
wire g17015;
wire g24269;
wire II18590;
wire II18710;
wire g29814;
wire g4369;
wire g16842;
wire g16643;
wire II21160;
wire g28915;
wire g20694;
wire g19521;
wire g22516;
wire g29989;
wire g29967;
wire g24317;
wire II28100;
wire g19984;
wire g7888;
wire g14177;
wire II13956;
wire II37781;
wire II31637;
wire g18166;
wire g30549;
wire g11683;
wire II35723;
wire g13933;
wire g8973;
wire g10883;
wire g4523;
wire II34863;
wire g16064;
wire II20299;
wire g29678;
wire II25222;
wire g16153;
wire g25472;
wire II38208;
wire g25698;
wire g10601;
wire g30067;
wire g11711;
wire g21301;
wire II16793;
wire II37617;
wire g21975;
wire g23179;
wire g7700;
wire g20735;
wire g11312;
wire II26401;
wire II22972;
wire g11516;
wire g16394;
wire g30597;
wire g29486;
wire g28317;
wire g7865;
wire g12461;
wire g4902;
wire II33837;
wire g4668;
wire g19596;
wire g19865;
wire g19708;
wire g16178;
wire g20400;
wire g24162;
wire g30695;
wire g8522;
wire II36939;
wire g11497;
wire II23923;
wire g22134;
wire g13863;
wire II40679;
wire II23123;
wire g19241;
wire II18184;
wire g9666;
wire g4281;
wire g9143;
wire g5685;
wire g4360;
wire g23232;
wire g22487;
wire g26335;
wire g9303;
wire g19109;
wire g4055;
wire g16299;
wire g19823;
wire g18245;
wire g15526;
wire g4754;
wire g29432;
wire g15411;
wire g9229;
wire g13354;
wire g15492;
wire g8230;
wire g15382;
wire g28768;
wire II25571;
wire g21802;
wire II36888;
wire g25844;
wire g9880;
wire g28133;
wire g10641;
wire II13538;
wire II29999;
wire g12119;
wire g28011;
wire g28332;
wire g20463;
wire g10909;
wire g13289;
wire g26151;
wire g12042;
wire g19556;
wire g21401;
wire g12597;
wire II40565;
wire g6042;
wire g29889;
wire II38128;
wire II24171;
wire g29519;
wire g19928;
wire II25264;
wire g7858;
wire g23258;
wire g23169;
wire g12881;
wire g21255;
wire II35814;
wire II30844;
wire II40251;
wire g13519;
wire II33232;
wire g27376;
wire g25392;
wire g12295;
wire g27501;
wire II30056;
wire g13029;
wire g26040;
wire gbuf32;
wire gbuf48;
wire g16476;
wire II32112;
wire II16664;
wire g9730;
wire g10623;
wire II23424;
wire g7739;
wire g16480;
wire II37880;
wire g18483;
wire II29418;
wire g5692;
wire II22575;
wire II29197;
wire g18088;
wire gbuf28;
wire II30547;
wire II16279;
wire II38080;
wire II31703;
wire g11243;
wire g11704;
wire II16131;
wire g18857;
wire g10412;
wire g21757;
wire II34086;
wire gbuf87;
wire II22618;
wire g5755;
wire II22611;
wire g21893;
wire g15887;
wire g14711;
wire g22150;
wire g16046;
wire g20296;
wire g28998;
wire g28699;
wire g5266;
wire g30763;
wire II39398;
wire II39674;
wire g21004;
wire g11846;
wire II20541;
wire g14991;
wire g23058;
wire g12471;
wire g16053;
wire II27029;
wire II14990;
wire II15602;
wire II14587;
wire II23527;
wire g11252;
wire g10573;
wire II24362;
wire g18307;
wire g24504;
wire II34096;
wire g26878;
wire II17235;
wire II34220;
wire g27695;
wire II27749;
wire g15435;
wire II35791;
wire g22227;
wire gbuf154;
wire g23438;
wire g4942;
wire g30671;
wire II36371;
wire II29939;
wire g3461;
wire g13452;
wire g29467;
wire g20892;
wire g20310;
wire II13143;
wire g27771;
wire II39026;
wire g25729;
wire g30770;
wire II22414;
wire II15350;
wire g17419;
wire g12657;
wire II25365;
wire g24036;
wire g27364;
wire g25173;
wire II37871;
wire g25523;
wire g20452;
wire g16676;
wire g28685;
wire g25761;
wire g9787;
wire gbuf140;
wire g22761;
wire g13317;
wire g13121;
wire g29298;
wire g23248;
wire g14347;
wire g13035;
wire g21781;
wire g28512;
wire g5394;
wire gbuf59;
wire g19727;
wire g15074;
wire g4955;
wire II29468;
wire II14865;
wire g26193;
wire g24057;
wire g15678;
wire g4301;
wire g26505;
wire g12821;
wire II34277;
wire g28232;
wire II24647;
wire II36072;
wire g21874;
wire g26347;
wire g10915;
wire II37752;
wire II21252;
wire g14546;
wire g10388;
wire g21670;
wire g24487;
wire II17756;
wire g15588;
wire g5728;
wire g5320;
wire g28079;
wire g19945;
wire II29579;
wire g16418;
wire g11567;
wire g18930;
wire g26852;
wire II33347;
wire II28178;
wire II19997;
wire II26612;
wire II18990;
wire g24856;
wire II37146;
wire II39237;
wire g23678;
wire II40495;
wire g4836;
wire g30678;
wire g8770;
wire II35394;
wire g26182;
wire g19012;
wire II23591;
wire g28152;
wire g16599;
wire g24757;
wire II30377;
wire g24773;
wire g19768;
wire II33790;
wire g7910;
wire II22999;
wire g13907;
wire g16140;
wire g12543;
wire g20430;
wire g16414;
wire g20411;
wire II20417;
wire g24574;
wire g23896;
wire g19194;
wire g19577;
wire g15609;
wire g20040;
wire g27464;
wire g15201;
wire g8726;
wire g8093;
wire g25714;
wire g5717;
wire g18222;
wire g29474;
wire II26661;
wire g11888;
wire g29570;
wire g24449;
wire g4139;
wire II32347;
wire II18323;
wire II40450;
wire g12363;
wire g11341;
wire g7580;
wire g17218;
wire g30297;
wire II36667;
wire g23038;
wire g19482;
wire II23008;
wire g23414;
wire g24491;
wire g23823;
wire g12513;
wire g17576;
wire g22597;
wire II31583;
wire g18815;
wire g25246;
wire g5957;
wire gbuf169;
wire g9423;
wire II27092;
wire g11417;
wire II17789;
wire g7333;
wire II29354;
wire g26671;
wire g11294;
wire g30988;
wire g10767;
wire g8792;
wire g7837;
wire g6161;
wire II40614;
wire II33501;
wire g30101;
wire g10796;
wire g11920;
wire g22629;
wire g24964;
wire g25212;
wire g23477;
wire g4976;
wire g13133;
wire gbuf202;
wire g7642;
wire g20966;
wire g27391;
wire g25278;
wire g10848;
wire g23273;
wire g22995;
wire II16206;
wire g29760;
wire II38613;
wire g15425;
wire g25404;
wire II19901;
wire g25631;
wire g19653;
wire g25457;
wire g19456;
wire II24624;
wire g23237;
wire II29506;
wire g12755;
wire g13352;
wire g18212;
wire g28971;
wire g26771;
wire g22130;
wire g29187;
wire g17926;
wire g21028;
wire g8028;
wire g5113;
wire g27897;
wire g13260;
wire g15544;
wire g15596;
wire g26249;
wire g26705;
wire g19657;
wire g29576;
wire II31053;
wire II16741;
wire g21990;
wire II41117;
wire g24748;
wire II14056;
wire g16859;
wire g28227;
wire g22263;
wire g30289;
wire g29285;
wire g22172;
wire g8153;
wire g20045;
wire g23132;
wire g22049;
wire II33268;
wire II40161;
wire g29158;
wire II33819;
wire II36972;
wire g21210;
wire II16325;
wire g30754;
wire g26550;
wire g29167;
wire II27766;
wire II29313;
wire g30591;
wire g27599;
wire g20349;
wire g20001;
wire g27238;
wire g30669;
wire II29058;
wire g25422;
wire g15284;
wire g23239;
wire g8538;
wire g26351;
wire II16857;
wire g25076;
wire II16482;
wire g19200;
wire g29343;
wire g12219;
wire g20884;
wire g16430;
wire g29708;
wire g22097;
wire g13426;
wire II26846;
wire g17490;
wire II36081;
wire g23435;
wire g7478;
wire g29039;
wire II31302;
wire g25944;
wire II14191;
wire II27658;
wire g24660;
wire g23151;
wire g27110;
wire g18678;
wire II20379;
wire g29307;
wire g10567;
wire II39926;
wire II25219;
wire g29275;
wire g10116;
wire g23319;
wire II30224;
wire g23470;
wire g22242;
wire g21336;
wire II16850;
wire g30970;
wire g30712;
wire II23287;
wire g28063;
wire g23014;
wire g13244;
wire g24555;
wire g16103;
wire g17754;
wire g22826;
wire II39828;
wire g15308;
wire II15562;
wire g21391;
wire g10093;
wire g5911;
wire II24566;
wire g27158;
wire g19281;
wire g26575;
wire g12959;
wire II25402;
wire g23938;
wire g24885;
wire g4089;
wire II29569;
wire g13224;
wire II29043;
wire II39690;
wire g10590;
wire II26558;
wire g13833;
wire g11303;
wire II35020;
wire II29924;
wire g17746;
wire g5404;
wire II40447;
wire II31517;
wire g22872;
wire g22062;
wire II39080;
wire g13099;
wire g20361;
wire g12425;
wire g25051;
wire II37035;
wire g15566;
wire g15423;
wire g8285;
wire g24152;
wire II33448;
wire g11003;
wire g25410;
wire g21742;
wire g30533;
wire II25374;
wire g12791;
wire g15357;
wire g22418;
wire g19022;
wire g18918;
wire II40670;
wire g30339;
wire g29338;
wire II37014;
wire g5844;
wire II19736;
wire g26060;
wire gbuf80;
wire g25882;
wire g28993;
wire g22113;
wire II38812;
wire g17395;
wire g7015;
wire g3254;
wire g21765;
wire g27066;
wire II19711;
wire II23057;
wire g18651;
wire II17804;
wire II40059;
wire g8351;
wire g19743;
wire g17919;
wire g29068;
wire II33822;
wire g28672;
wire II21586;
wire g26008;
wire g21147;
wire g24071;
wire g22991;
wire g26382;
wire II18554;
wire g21912;
wire II39391;
wire II36337;
wire g24534;
wire g12001;
wire g4693;
wire g10198;
wire g11082;
wire g30600;
wire g28031;
wire II17527;
wire g15225;
wire g17697;
wire g23785;
wire g18205;
wire g23418;
wire g11553;
wire g18463;
wire g13239;
wire g27313;
wire g29621;
wire II15299;
wire g27472;
wire II33636;
wire g19223;
wire II32266;
wire g27176;
wire II24718;
wire g27810;
wire II27221;
wire g25943;
wire II23199;
wire g5167;
wire g19094;
wire g30664;
wire g13419;
wire II14238;
wire g16487;
wire II29392;
wire II29151;
wire g17130;
wire g18913;
wire g24000;
wire g25273;
wire g24516;
wire II33627;
wire II32401;
wire g3251;
wire g29645;
wire g21228;
wire g27179;
wire g23566;
wire II34824;
wire g13414;
wire g28427;
wire g10445;
wire II38056;
wire g30237;
wire g5898;
wire II25528;
wire g10285;
wire II28767;
wire g16110;
wire II29262;
wire g23820;
wire g17893;
wire g6304;
wire g10859;
wire II31014;
wire g17028;
wire g20107;
wire g12945;
wire g30654;
wire II21277;
wire g24046;
wire g12951;
wire g29978;
wire II31270;
wire II27422;
wire g20584;
wire g22674;
wire II24213;
wire II30826;
wire II30651;
wire g25271;
wire g17842;
wire g24250;
wire g23973;
wire g23747;
wire g20112;
wire g27755;
wire II39086;
wire g18772;
wire g16171;
wire g26399;
wire II35744;
wire II16939;
wire g21438;
wire g29697;
wire g21039;
wire g25724;
wire II18169;
wire II36769;
wire g29920;
wire g5015;
wire g21866;
wire g12521;
wire g21606;
wire g10931;
wire II23942;
wire gbuf132;
wire g13496;
wire g5640;
wire g20500;
wire g14618;
wire II33577;
wire II32934;
wire g13143;
wire II22925;
wire g29476;
wire g15322;
wire gbuf149;
wire II25096;
wire g23719;
wire g11747;
wire II39906;
wire g23260;
wire II36975;
wire II40134;
wire II35022;
wire II30308;
wire g25780;
wire g20545;
wire g15623;
wire g24228;
wire g30769;
wire g9161;
wire II39463;
wire g27734;
wire g28368;
wire g4862;
wire II38692;
wire g12129;
wire g8650;
wire g22222;
wire g25120;
wire II31159;
wire g27187;
wire II15574;
wire g18890;
wire II21259;
wire g28445;
wire gbuf58;
wire g15878;
wire g13100;
wire II30480;
wire g28823;
wire II13677;
wire II25839;
wire g8811;
wire g26653;
wire g21252;
wire II22632;
wire g30557;
wire II19615;
wire II32210;
wire g23734;
wire g4869;
wire g25552;
wire g18079;
wire g10966;
wire g30381;
wire II40922;
wire g23554;
wire g4165;
wire g10211;
wire g21061;
wire II15238;
wire g9733;
wire g13943;
wire g18780;
wire g19690;
wire g20825;
wire g11912;
wire g23906;
wire g15176;
wire g4860;
wire g3305;
wire g19632;
wire g27486;
wire g11985;
wire II26491;
wire II36636;
wire g13188;
wire g10409;
wire g10404;
wire g28618;
wire g6030;
wire g24836;
wire g15704;
wire g19906;
wire g10398;
wire g7852;
wire g5000;
wire g4260;
wire II39803;
wire II20667;
wire g24369;
wire g18841;
wire II34967;
wire g3866;
wire g15261;
wire g13094;
wire II28896;
wire g13335;
wire g25350;
wire g8933;
wire g30719;
wire II40182;
wire g8705;
wire II34074;
wire II16450;
wire g16491;
wire g20630;
wire II24667;
wire g21619;
wire g20222;
wire g26669;
wire g25222;
wire g17168;
wire II31035;
wire II16341;
wire g5301;
wire g22287;
wire II38091;
wire II33673;
wire II37497;
wire g19135;
wire II20506;
wire II31553;
wire g23672;
wire g5596;
wire II23775;
wire g25499;
wire g16390;
wire g14502;
wire g11903;
wire g3493;
wire g27738;
wire g17554;
wire II30140;
wire II34848;
wire II20607;
wire II18037;
wire g5933;
wire g9954;
wire II30110;
wire II28330;
wire g26051;
wire II27405;
wire g26268;
wire II34704;
wire g13655;
wire II31037;
wire g27291;
wire g9632;
wire II39641;
wire g4224;
wire g17461;
wire g12009;
wire g13384;
wire II38085;
wire g4143;
wire II35479;
wire g22190;
wire g17354;
wire g23517;
wire g17499;
wire g24065;
wire g26279;
wire g16824;
wire g27699;
wire II27101;
wire g12749;
wire g13904;
wire g22156;
wire g29092;
wire g25506;
wire g26759;
wire II31091;
wire g23298;
wire II25830;
wire g21772;
wire g8506;
wire g9910;
wire g22331;
wire g10130;
wire II15463;
wire II35007;
wire g24345;
wire g29682;
wire II15317;
wire g21612;
wire g4674;
wire g17137;
wire g24375;
wire g21481;
wire g4124;
wire g12944;
wire g21739;
wire II23412;
wire g26715;
wire II38238;
wire g6104;
wire g19348;
wire II40531;
wire g22584;
wire g27426;
wire g26830;
wire g10788;
wire g6053;
wire II30952;
wire g17479;
wire II15184;
wire g28847;
wire g6043;
wire g22280;
wire g25230;
wire II28800;
wire II18503;
wire g21790;
wire II25771;
wire g24907;
wire g24924;
wire g10322;
wire II21491;
wire g11560;
wire g27081;
wire II39047;
wire g28293;
wire g16034;
wire g19050;
wire II33431;
wire g24401;
wire g24900;
wire II36468;
wire g29304;
wire II23364;
wire g23802;
wire II38345;
wire II17857;
wire g19089;
wire II35044;
wire g11861;
wire g30222;
wire g26494;
wire g10933;
wire II20743;
wire g29391;
wire II21942;
wire g27722;
wire II18113;
wire g7542;
wire g12552;
wire g9952;
wire g28210;
wire g24319;
wire g17875;
wire II35099;
wire g17047;
wire II28057;
wire II14834;
wire g11641;
wire g11814;
wire g21690;
wire g5938;
wire II40946;
wire g23982;
wire g14123;
wire II34752;
wire g30068;
wire g21794;
wire g23139;
wire g13571;
wire g5088;
wire II32976;
wire g5828;
wire II29323;
wire g4438;
wire II37101;
wire II23788;
wire g8408;
wire g16036;
wire g27180;
wire g20924;
wire II32928;
wire g29016;
wire g29314;
wire g27908;
wire g24758;
wire g13359;
wire II20467;
wire II32697;
wire II39635;
wire g8870;
wire g12305;
wire II21905;
wire g23837;
wire II32907;
wire g20188;
wire II24049;
wire II29903;
wire g30092;
wire II30901;
wire g25590;
wire g22275;
wire g13160;
wire g17145;
wire II34244;
wire II39942;
wire g8491;
wire g16758;
wire g28167;
wire II39540;
wire II33852;
wire g19231;
wire g26811;
wire II29165;
wire g21747;
wire g26631;
wire g22990;
wire II15654;
wire g13467;
wire g30473;
wire g6079;
wire g29783;
wire II16053;
wire g19575;
wire II28969;
wire g22267;
wire II39821;
wire II14942;
wire II27074;
wire g30826;
wire g15037;
wire g27336;
wire g12840;
wire II18311;
wire g18004;
wire g20941;
wire g30792;
wire g10704;
wire g15869;
wire g23111;
wire g8498;
wire g30304;
wire II37793;
wire II39005;
wire g11025;
wire g24351;
wire II25231;
wire g11535;
wire g15999;
wire II37056;
wire II31226;
wire g28240;
wire g13191;
wire g24183;
wire II32333;
wire g13107;
wire II16037;
wire g11726;
wire g26280;
wire II19883;
wire g21528;
wire g18807;
wire g12409;
wire II23292;
wire g24435;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2814 <= 0;
  else
    g2814 <= g16475;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2817 <= 0;
  else
    g2817 <= g20571;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2933 <= 0;
  else
    g2933 <= g20588;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2950 <= 0;
  else
    g2950 <= g21951;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2883 <= 0;
  else
    g2883 <= g23315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2888 <= 0;
  else
    g2888 <= g24423;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2896 <= 0;
  else
    g2896 <= g25175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2892 <= 0;
  else
    g2892 <= g26019;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2903 <= 0;
  else
    g2903 <= g26747;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2900 <= 0;
  else
    g2900 <= g27237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2908 <= 0;
  else
    g2908 <= g27715;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2912 <= 0;
  else
    g2912 <= g24424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2917 <= 0;
  else
    g2917 <= g25174;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2924 <= 0;
  else
    g2924 <= g26020;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2920 <= 0;
  else
    g2920 <= g26746;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2984 <= 0;
  else
    g2984 <= g19061;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2985 <= 0;
  else
    g2985 <= g19060;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2930 <= 0;
  else
    g2930 <= g19062;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2929 <= 0;
  else
    g2929 <= gbuf1;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2879 <= 0;
  else
    g2879 <= g16494;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2934 <= 0;
  else
    g2934 <= g16476;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2935 <= 0;
  else
    g2935 <= g16477;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2938 <= 0;
  else
    g2938 <= g16478;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2941 <= 0;
  else
    g2941 <= g16479;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2944 <= 0;
  else
    g2944 <= g16480;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2947 <= 0;
  else
    g2947 <= g16481;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2953 <= 0;
  else
    g2953 <= g16482;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2956 <= 0;
  else
    g2956 <= g16483;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2959 <= 0;
  else
    g2959 <= g16484;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2962 <= 0;
  else
    g2962 <= g16485;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2963 <= 0;
  else
    g2963 <= g16486;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2966 <= 0;
  else
    g2966 <= g16487;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2969 <= 0;
  else
    g2969 <= g16488;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2972 <= 0;
  else
    g2972 <= g16489;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2975 <= 0;
  else
    g2975 <= g16490;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2978 <= 0;
  else
    g2978 <= g16491;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2981 <= 0;
  else
    g2981 <= g16492;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2874 <= 0;
  else
    g2874 <= g16493;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1506 <= 0;
  else
    g1506 <= g20572;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1501 <= 0;
  else
    g1501 <= g20573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1496 <= 0;
  else
    g1496 <= g20574;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1491 <= 0;
  else
    g1491 <= g20575;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1486 <= 0;
  else
    g1486 <= g20576;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1481 <= 0;
  else
    g1481 <= g20577;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1476 <= 0;
  else
    g1476 <= g20578;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1471 <= 0;
  else
    g1471 <= g20579;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2877 <= 0;
  else
    g2877 <= g23313;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2861 <= 0;
  else
    g2861 <= g21960;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g813 <= 0;
  else
    g813 <= gbuf2;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2864 <= 0;
  else
    g2864 <= g21961;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g809 <= 0;
  else
    g809 <= gbuf3;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2867 <= 0;
  else
    g2867 <= g21962;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g805 <= 0;
  else
    g805 <= gbuf4;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2870 <= 0;
  else
    g2870 <= g21963;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g801 <= 0;
  else
    g801 <= gbuf5;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2818 <= 0;
  else
    g2818 <= g21947;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g797 <= 0;
  else
    g797 <= gbuf6;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2821 <= 0;
  else
    g2821 <= g21948;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g793 <= 0;
  else
    g793 <= gbuf7;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2824 <= 0;
  else
    g2824 <= g21949;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g789 <= 0;
  else
    g789 <= gbuf8;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2827 <= 0;
  else
    g2827 <= g21950;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g785 <= 0;
  else
    g785 <= gbuf9;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2830 <= 0;
  else
    g2830 <= g23312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2873 <= 0;
  else
    g2873 <= gbuf10;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2833 <= 0;
  else
    g2833 <= g21952;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g125 <= 0;
  else
    g125 <= gbuf11;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2836 <= 0;
  else
    g2836 <= g21953;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g121 <= 0;
  else
    g121 <= gbuf12;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2839 <= 0;
  else
    g2839 <= g21954;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g117 <= 0;
  else
    g117 <= gbuf13;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2842 <= 0;
  else
    g2842 <= g21955;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g113 <= 0;
  else
    g113 <= gbuf14;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2845 <= 0;
  else
    g2845 <= g21956;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g109 <= 0;
  else
    g109 <= gbuf15;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2848 <= 0;
  else
    g2848 <= g21957;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g105 <= 0;
  else
    g105 <= gbuf16;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2851 <= 0;
  else
    g2851 <= g21958;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g101 <= 0;
  else
    g101 <= gbuf17;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2854 <= 0;
  else
    g2854 <= g21959;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g97 <= 0;
  else
    g97 <= gbuf18;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2858 <= 0;
  else
    g2858 <= g23316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2857 <= 0;
  else
    g2857 <= gbuf19;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2200 <= 0;
  else
    g2200 <= g20587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2195 <= 0;
  else
    g2195 <= g20585;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2190 <= 0;
  else
    g2190 <= g20586;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2185 <= 0;
  else
    g2185 <= g20584;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2180 <= 0;
  else
    g2180 <= g20583;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2175 <= 0;
  else
    g2175 <= g20582;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2170 <= 0;
  else
    g2170 <= g20581;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2165 <= 0;
  else
    g2165 <= g20580;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2878 <= 0;
  else
    g2878 <= g23314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3129 <= 0;
  else
    g3129 <= g13475;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3117 <= 0;
  else
    g3117 <= gbuf20;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3109 <= 0;
  else
    g3109 <= gbuf21;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3210 <= 0;
  else
    g3210 <= g20630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3211 <= 0;
  else
    g3211 <= g20631;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3084 <= 0;
  else
    g3084 <= g20632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3085 <= 0;
  else
    g3085 <= g20609;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3086 <= 0;
  else
    g3086 <= g20610;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3087 <= 0;
  else
    g3087 <= g20611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3091 <= 0;
  else
    g3091 <= g20612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3092 <= 0;
  else
    g3092 <= g20613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3093 <= 0;
  else
    g3093 <= g20614;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3094 <= 0;
  else
    g3094 <= g20615;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3095 <= 0;
  else
    g3095 <= g20616;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3096 <= 0;
  else
    g3096 <= g20617;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3097 <= 0;
  else
    g3097 <= g26751;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3098 <= 0;
  else
    g3098 <= g26752;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3099 <= 0;
  else
    g3099 <= g26753;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3100 <= 0;
  else
    g3100 <= g29163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3101 <= 0;
  else
    g3101 <= g29164;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3102 <= 0;
  else
    g3102 <= g29165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3103 <= 0;
  else
    g3103 <= g30120;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3104 <= 0;
  else
    g3104 <= g30121;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3105 <= 0;
  else
    g3105 <= g30122;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3106 <= 0;
  else
    g3106 <= g30941;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3107 <= 0;
  else
    g3107 <= g30942;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3108 <= 0;
  else
    g3108 <= g30943;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3155 <= 0;
  else
    g3155 <= g20618;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3158 <= 0;
  else
    g3158 <= g20619;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3161 <= 0;
  else
    g3161 <= g20620;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3164 <= 0;
  else
    g3164 <= g20621;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3167 <= 0;
  else
    g3167 <= g20622;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3170 <= 0;
  else
    g3170 <= g20623;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3173 <= 0;
  else
    g3173 <= g20624;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3176 <= 0;
  else
    g3176 <= g20625;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3179 <= 0;
  else
    g3179 <= g20626;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3182 <= 0;
  else
    g3182 <= g20627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3185 <= 0;
  else
    g3185 <= g20628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3088 <= 0;
  else
    g3088 <= g20629;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3191 <= 0;
  else
    g3191 <= g27717;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3194 <= 0;
  else
    g3194 <= g28316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3197 <= 0;
  else
    g3197 <= g28317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3198 <= 0;
  else
    g3198 <= g28318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3201 <= 0;
  else
    g3201 <= g28704;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3204 <= 0;
  else
    g3204 <= g28705;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3207 <= 0;
  else
    g3207 <= g28706;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3188 <= 0;
  else
    g3188 <= g29463;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3133 <= 0;
  else
    g3133 <= g29656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3132 <= 0;
  else
    g3132 <= g28698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3128 <= 0;
  else
    g3128 <= g29166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3127 <= 0;
  else
    g3127 <= g28697;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3126 <= 0;
  else
    g3126 <= g28315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3125 <= 0;
  else
    g3125 <= g28696;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3124 <= 0;
  else
    g3124 <= g28314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3123 <= 0;
  else
    g3123 <= g28313;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3120 <= 0;
  else
    g3120 <= g28695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3114 <= 0;
  else
    g3114 <= g28694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3113 <= 0;
  else
    g3113 <= g28693;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3112 <= 0;
  else
    g3112 <= g28312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3110 <= 0;
  else
    g3110 <= g28311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3111 <= 0;
  else
    g3111 <= g28310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3139 <= 0;
  else
    g3139 <= g29461;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3136 <= 0;
  else
    g3136 <= g28701;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3134 <= 0;
  else
    g3134 <= g28700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3135 <= 0;
  else
    g3135 <= g28699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3151 <= 0;
  else
    g3151 <= g29462;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3142 <= 0;
  else
    g3142 <= g28703;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3147 <= 0;
  else
    g3147 <= g28702;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g185 <= 0;
  else
    g185 <= g29657;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g138 <= 0;
  else
    g138 <= g13405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g135 <= 0;
  else
    g135 <= gbuf22;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g165 <= 0;
  else
    g165 <= gbuf23;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g130 <= 0;
  else
    g130 <= g24259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g131 <= 0;
  else
    g131 <= g24260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g129 <= 0;
  else
    g129 <= g24261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g133 <= 0;
  else
    g133 <= g24262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g134 <= 0;
  else
    g134 <= g24263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g132 <= 0;
  else
    g132 <= g24264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g142 <= 0;
  else
    g142 <= g24265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g143 <= 0;
  else
    g143 <= g24266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g141 <= 0;
  else
    g141 <= g24267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g145 <= 0;
  else
    g145 <= g24268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g146 <= 0;
  else
    g146 <= g24269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g144 <= 0;
  else
    g144 <= g24270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g148 <= 0;
  else
    g148 <= g24271;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g149 <= 0;
  else
    g149 <= g24272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g147 <= 0;
  else
    g147 <= g24273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g151 <= 0;
  else
    g151 <= g24274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g152 <= 0;
  else
    g152 <= g24275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g150 <= 0;
  else
    g150 <= g24276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g154 <= 0;
  else
    g154 <= g24277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g155 <= 0;
  else
    g155 <= g24278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g153 <= 0;
  else
    g153 <= g24279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g157 <= 0;
  else
    g157 <= g24280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g158 <= 0;
  else
    g158 <= g24281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g156 <= 0;
  else
    g156 <= g24282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g160 <= 0;
  else
    g160 <= g24283;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g161 <= 0;
  else
    g161 <= g24284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g159 <= 0;
  else
    g159 <= g24285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g163 <= 0;
  else
    g163 <= g24286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g164 <= 0;
  else
    g164 <= g24287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g162 <= 0;
  else
    g162 <= g24288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g169 <= 0;
  else
    g169 <= g26679;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g170 <= 0;
  else
    g170 <= g26680;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g168 <= 0;
  else
    g168 <= g26681;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g172 <= 0;
  else
    g172 <= g26682;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g173 <= 0;
  else
    g173 <= g26683;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g171 <= 0;
  else
    g171 <= g26684;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g175 <= 0;
  else
    g175 <= g26685;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g176 <= 0;
  else
    g176 <= g26686;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g174 <= 0;
  else
    g174 <= g26687;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g178 <= 0;
  else
    g178 <= g26688;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g179 <= 0;
  else
    g179 <= g26689;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g177 <= 0;
  else
    g177 <= g26690;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g186 <= 0;
  else
    g186 <= g30506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g189 <= 0;
  else
    g189 <= g30507;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g192 <= 0;
  else
    g192 <= g30508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g231 <= 0;
  else
    g231 <= g30842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g234 <= 0;
  else
    g234 <= g30843;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g237 <= 0;
  else
    g237 <= g30844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g195 <= 0;
  else
    g195 <= g30836;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g198 <= 0;
  else
    g198 <= g30837;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g201 <= 0;
  else
    g201 <= g30838;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g240 <= 0;
  else
    g240 <= g30845;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g243 <= 0;
  else
    g243 <= g30846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g246 <= 0;
  else
    g246 <= g30847;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g204 <= 0;
  else
    g204 <= g30509;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g207 <= 0;
  else
    g207 <= g30510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g210 <= 0;
  else
    g210 <= g30511;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g249 <= 0;
  else
    g249 <= g30515;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g252 <= 0;
  else
    g252 <= g30516;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g255 <= 0;
  else
    g255 <= g30517;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g213 <= 0;
  else
    g213 <= g30512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g216 <= 0;
  else
    g216 <= g30513;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g219 <= 0;
  else
    g219 <= g30514;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g258 <= 0;
  else
    g258 <= g30518;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g261 <= 0;
  else
    g261 <= g30519;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g264 <= 0;
  else
    g264 <= g30520;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g222 <= 0;
  else
    g222 <= g30839;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g225 <= 0;
  else
    g225 <= g30840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g228 <= 0;
  else
    g228 <= g30841;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g267 <= 0;
  else
    g267 <= g30848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g270 <= 0;
  else
    g270 <= g30849;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g273 <= 0;
  else
    g273 <= g30850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g92 <= 0;
  else
    g92 <= g25983;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g88 <= 0;
  else
    g88 <= g26678;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g83 <= 0;
  else
    g83 <= g27189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g79 <= 0;
  else
    g79 <= g27683;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g74 <= 0;
  else
    g74 <= g28206;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g70 <= 0;
  else
    g70 <= g28673;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g65 <= 0;
  else
    g65 <= g29131;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g61 <= 0;
  else
    g61 <= g29413;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g56 <= 0;
  else
    g56 <= g29627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g52 <= 0;
  else
    g52 <= g29794;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g180 <= 0;
  else
    g180 <= g20555;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g182 <= 0;
  else
    g182 <= gbuf24;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g181 <= 0;
  else
    g181 <= gbuf25;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g276 <= 0;
  else
    g276 <= g13406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g405 <= 0;
  else
    g405 <= gbuf26;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g401 <= 0;
  else
    g401 <= gbuf27;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g309 <= 0;
  else
    g309 <= g11496;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g354 <= 0;
  else
    g354 <= g28207;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g343 <= 0;
  else
    g343 <= g28208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g346 <= 0;
  else
    g346 <= g28209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g369 <= 0;
  else
    g369 <= g28210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g358 <= 0;
  else
    g358 <= g28211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g361 <= 0;
  else
    g361 <= g28212;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g384 <= 0;
  else
    g384 <= g28213;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g373 <= 0;
  else
    g373 <= g28214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g376 <= 0;
  else
    g376 <= g28215;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g398 <= 0;
  else
    g398 <= g28216;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g388 <= 0;
  else
    g388 <= g28217;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g391 <= 0;
  else
    g391 <= g28218;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g408 <= 0;
  else
    g408 <= g29414;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g411 <= 0;
  else
    g411 <= g29415;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g414 <= 0;
  else
    g414 <= g29416;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g417 <= 0;
  else
    g417 <= g29631;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g420 <= 0;
  else
    g420 <= g29632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g423 <= 0;
  else
    g423 <= g29633;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g427 <= 0;
  else
    g427 <= g29417;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g428 <= 0;
  else
    g428 <= g29418;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g426 <= 0;
  else
    g426 <= g29419;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g429 <= 0;
  else
    g429 <= g27684;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g432 <= 0;
  else
    g432 <= g27685;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g435 <= 0;
  else
    g435 <= g27686;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g438 <= 0;
  else
    g438 <= g27687;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g441 <= 0;
  else
    g441 <= g27688;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g444 <= 0;
  else
    g444 <= g27689;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g448 <= 0;
  else
    g448 <= g28674;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g449 <= 0;
  else
    g449 <= g28675;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g447 <= 0;
  else
    g447 <= g28676;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g312 <= 0;
  else
    g312 <= g29795;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g313 <= 0;
  else
    g313 <= g29796;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g314 <= 0;
  else
    g314 <= g29797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g315 <= 0;
  else
    g315 <= g30851;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g316 <= 0;
  else
    g316 <= g30852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g317 <= 0;
  else
    g317 <= g30853;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g318 <= 0;
  else
    g318 <= g30710;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g319 <= 0;
  else
    g319 <= g30711;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g320 <= 0;
  else
    g320 <= g30712;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g322 <= 0;
  else
    g322 <= g29628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g323 <= 0;
  else
    g323 <= g29629;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g321 <= 0;
  else
    g321 <= g29630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g403 <= 0;
  else
    g403 <= g27191;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g404 <= 0;
  else
    g404 <= g27192;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g402 <= 0;
  else
    g402 <= g27193;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g450 <= 0;
  else
    g450 <= g11509;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g451 <= 0;
  else
    g451 <= gbuf28;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g452 <= 0;
  else
    g452 <= g11510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g453 <= 0;
  else
    g453 <= gbuf29;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g454 <= 0;
  else
    g454 <= g11511;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g279 <= 0;
  else
    g279 <= gbuf30;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g280 <= 0;
  else
    g280 <= g11491;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g281 <= 0;
  else
    g281 <= gbuf31;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g282 <= 0;
  else
    g282 <= g11492;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g283 <= 0;
  else
    g283 <= gbuf32;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g284 <= 0;
  else
    g284 <= g11493;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g285 <= 0;
  else
    g285 <= gbuf33;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g286 <= 0;
  else
    g286 <= g11494;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g287 <= 0;
  else
    g287 <= gbuf34;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g288 <= 0;
  else
    g288 <= g11495;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g289 <= 0;
  else
    g289 <= gbuf35;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g290 <= 0;
  else
    g290 <= g13407;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g291 <= 0;
  else
    g291 <= gbuf36;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g299 <= 0;
  else
    g299 <= g19012;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g305 <= 0;
  else
    g305 <= g23148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g308 <= 0;
  else
    g308 <= g23149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g297 <= 0;
  else
    g297 <= g23150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g296 <= 0;
  else
    g296 <= g23151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g295 <= 0;
  else
    g295 <= g23152;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g294 <= 0;
  else
    g294 <= g23153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g304 <= 0;
  else
    g304 <= g19016;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g303 <= 0;
  else
    g303 <= g19015;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g302 <= 0;
  else
    g302 <= g19014;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g301 <= 0;
  else
    g301 <= g19013;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g300 <= 0;
  else
    g300 <= g25130;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g298 <= 0;
  else
    g298 <= g27190;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g342 <= 0;
  else
    g342 <= g11497;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g349 <= 0;
  else
    g349 <= gbuf37;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g350 <= 0;
  else
    g350 <= g11498;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g351 <= 0;
  else
    g351 <= gbuf38;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g352 <= 0;
  else
    g352 <= g11499;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g353 <= 0;
  else
    g353 <= gbuf39;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g357 <= 0;
  else
    g357 <= g11500;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g364 <= 0;
  else
    g364 <= gbuf40;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g365 <= 0;
  else
    g365 <= g11501;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g366 <= 0;
  else
    g366 <= gbuf41;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g367 <= 0;
  else
    g367 <= g11502;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g368 <= 0;
  else
    g368 <= gbuf42;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g372 <= 0;
  else
    g372 <= g11503;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g379 <= 0;
  else
    g379 <= gbuf43;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g380 <= 0;
  else
    g380 <= g11504;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g381 <= 0;
  else
    g381 <= gbuf44;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g382 <= 0;
  else
    g382 <= g11505;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g383 <= 0;
  else
    g383 <= gbuf45;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g387 <= 0;
  else
    g387 <= g11506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g394 <= 0;
  else
    g394 <= gbuf46;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g395 <= 0;
  else
    g395 <= g11507;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g396 <= 0;
  else
    g396 <= gbuf47;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g397 <= 0;
  else
    g397 <= g11508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g324 <= 0;
  else
    g324 <= gbuf48;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g325 <= 0;
  else
    g325 <= g13408;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g331 <= 0;
  else
    g331 <= gbuf49;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g337 <= 0;
  else
    g337 <= gbuf50;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g545 <= 0;
  else
    g545 <= g13419;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g551 <= 0;
  else
    g551 <= gbuf51;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g550 <= 0;
  else
    g550 <= gbuf52;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g554 <= 0;
  else
    g554 <= g23160;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g557 <= 0;
  else
    g557 <= g20556;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g510 <= 0;
  else
    g510 <= g20557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g513 <= 0;
  else
    g513 <= g16467;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g523 <= 0;
  else
    g523 <= gbuf53;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g524 <= 0;
  else
    g524 <= gbuf54;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g564 <= 0;
  else
    g564 <= g11512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g569 <= 0;
  else
    g569 <= gbuf55;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g570 <= 0;
  else
    g570 <= g11515;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g571 <= 0;
  else
    g571 <= gbuf56;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g572 <= 0;
  else
    g572 <= g11516;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g573 <= 0;
  else
    g573 <= gbuf57;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g574 <= 0;
  else
    g574 <= g11517;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g565 <= 0;
  else
    g565 <= gbuf58;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g566 <= 0;
  else
    g566 <= g11513;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g567 <= 0;
  else
    g567 <= gbuf59;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g568 <= 0;
  else
    g568 <= g11514;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g489 <= 0;
  else
    g489 <= gbuf60;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g474 <= 0;
  else
    g474 <= g13409;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g481 <= 0;
  else
    g481 <= gbuf61;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g485 <= 0;
  else
    g485 <= gbuf62;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g486 <= 0;
  else
    g486 <= g24292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g487 <= 0;
  else
    g487 <= g24293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g488 <= 0;
  else
    g488 <= g24294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g455 <= 0;
  else
    g455 <= g25139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g458 <= 0;
  else
    g458 <= g25131;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g461 <= 0;
  else
    g461 <= g25132;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g477 <= 0;
  else
    g477 <= g25136;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g478 <= 0;
  else
    g478 <= g25137;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g479 <= 0;
  else
    g479 <= g25138;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g480 <= 0;
  else
    g480 <= g24289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g484 <= 0;
  else
    g484 <= g24290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g464 <= 0;
  else
    g464 <= g24291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g465 <= 0;
  else
    g465 <= g25133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g468 <= 0;
  else
    g468 <= g25134;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g471 <= 0;
  else
    g471 <= g25135;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g528 <= 0;
  else
    g528 <= g16468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g535 <= 0;
  else
    g535 <= gbuf63;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g542 <= 0;
  else
    g542 <= gbuf64;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g543 <= 0;
  else
    g543 <= g19021;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g544 <= 0;
  else
    g544 <= gbuf65;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g548 <= 0;
  else
    g548 <= g23159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g549 <= 0;
  else
    g549 <= g19022;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g499 <= 0;
  else
    g499 <= gbuf66;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g558 <= 0;
  else
    g558 <= g19023;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g559 <= 0;
  else
    g559 <= gbuf67;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g576 <= 0;
  else
    g576 <= g28219;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g577 <= 0;
  else
    g577 <= g28220;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g575 <= 0;
  else
    g575 <= g28221;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g579 <= 0;
  else
    g579 <= g28222;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g580 <= 0;
  else
    g580 <= g28223;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g578 <= 0;
  else
    g578 <= g28224;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g582 <= 0;
  else
    g582 <= g28225;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g583 <= 0;
  else
    g583 <= g28226;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g581 <= 0;
  else
    g581 <= g28227;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g585 <= 0;
  else
    g585 <= g28228;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g586 <= 0;
  else
    g586 <= g28229;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g584 <= 0;
  else
    g584 <= g28230;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g587 <= 0;
  else
    g587 <= g25985;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g590 <= 0;
  else
    g590 <= g25986;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g593 <= 0;
  else
    g593 <= g25987;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g596 <= 0;
  else
    g596 <= g25988;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g599 <= 0;
  else
    g599 <= g25989;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g602 <= 0;
  else
    g602 <= g25990;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g614 <= 0;
  else
    g614 <= g29135;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g617 <= 0;
  else
    g617 <= g29136;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g620 <= 0;
  else
    g620 <= g29137;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g605 <= 0;
  else
    g605 <= g29132;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g608 <= 0;
  else
    g608 <= g29133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g611 <= 0;
  else
    g611 <= g29134;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g490 <= 0;
  else
    g490 <= g27194;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g493 <= 0;
  else
    g493 <= g27195;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g496 <= 0;
  else
    g496 <= g27196;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g506 <= 0;
  else
    g506 <= g8284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g507 <= 0;
  else
    g507 <= g24295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g508 <= 0;
  else
    g508 <= g19017;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g509 <= 0;
  else
    g509 <= g19018;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g514 <= 0;
  else
    g514 <= g19019;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g515 <= 0;
  else
    g515 <= g19020;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g516 <= 0;
  else
    g516 <= g23158;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g517 <= 0;
  else
    g517 <= g23157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g518 <= 0;
  else
    g518 <= g23156;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g519 <= 0;
  else
    g519 <= g23155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g520 <= 0;
  else
    g520 <= g23154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g525 <= 0;
  else
    g525 <= gbuf68;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g529 <= 0;
  else
    g529 <= g13410;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g530 <= 0;
  else
    g530 <= g13411;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g531 <= 0;
  else
    g531 <= g13412;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g532 <= 0;
  else
    g532 <= g13413;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g533 <= 0;
  else
    g533 <= g13414;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g534 <= 0;
  else
    g534 <= g13415;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g536 <= 0;
  else
    g536 <= g13416;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g537 <= 0;
  else
    g537 <= g13417;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g538 <= 0;
  else
    g538 <= g25984;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g541 <= 0;
  else
    g541 <= g13418;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g623 <= 0;
  else
    g623 <= g13420;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g626 <= 0;
  else
    g626 <= gbuf69;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g629 <= 0;
  else
    g629 <= gbuf70;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g630 <= 0;
  else
    g630 <= g20558;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g659 <= 0;
  else
    g659 <= g21943;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g640 <= 0;
  else
    g640 <= g23161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g633 <= 0;
  else
    g633 <= g24296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g653 <= 0;
  else
    g653 <= g25140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g646 <= 0;
  else
    g646 <= g25991;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g660 <= 0;
  else
    g660 <= g26691;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g672 <= 0;
  else
    g672 <= g27197;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g666 <= 0;
  else
    g666 <= g27690;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g679 <= 0;
  else
    g679 <= g28231;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g686 <= 0;
  else
    g686 <= g28677;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g692 <= 0;
  else
    g692 <= g29138;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g699 <= 0;
  else
    g699 <= g23162;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g700 <= 0;
  else
    g700 <= g23163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g698 <= 0;
  else
    g698 <= g23164;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g702 <= 0;
  else
    g702 <= g23165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g703 <= 0;
  else
    g703 <= g23166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g701 <= 0;
  else
    g701 <= g23167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g705 <= 0;
  else
    g705 <= g23168;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g706 <= 0;
  else
    g706 <= g23169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g704 <= 0;
  else
    g704 <= g23170;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g708 <= 0;
  else
    g708 <= g23171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g709 <= 0;
  else
    g709 <= g23172;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g707 <= 0;
  else
    g707 <= g23173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g711 <= 0;
  else
    g711 <= g23174;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g712 <= 0;
  else
    g712 <= g23175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g710 <= 0;
  else
    g710 <= g23176;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g714 <= 0;
  else
    g714 <= g23177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g715 <= 0;
  else
    g715 <= g23178;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g713 <= 0;
  else
    g713 <= g23179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g717 <= 0;
  else
    g717 <= g23180;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g718 <= 0;
  else
    g718 <= g23181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g716 <= 0;
  else
    g716 <= g23182;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g720 <= 0;
  else
    g720 <= g23183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g721 <= 0;
  else
    g721 <= g23184;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g719 <= 0;
  else
    g719 <= g23185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g723 <= 0;
  else
    g723 <= g23186;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g724 <= 0;
  else
    g724 <= g23187;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g722 <= 0;
  else
    g722 <= g23188;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g726 <= 0;
  else
    g726 <= g23189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g727 <= 0;
  else
    g727 <= g23190;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g725 <= 0;
  else
    g725 <= g23191;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g729 <= 0;
  else
    g729 <= g23192;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g730 <= 0;
  else
    g730 <= g23193;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g728 <= 0;
  else
    g728 <= g23194;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g732 <= 0;
  else
    g732 <= g23195;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g733 <= 0;
  else
    g733 <= g23196;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g731 <= 0;
  else
    g731 <= g23197;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g735 <= 0;
  else
    g735 <= g26692;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g736 <= 0;
  else
    g736 <= g26693;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g734 <= 0;
  else
    g734 <= g26694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g738 <= 0;
  else
    g738 <= g24297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g739 <= 0;
  else
    g739 <= g24298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g737 <= 0;
  else
    g737 <= g24299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g826 <= 0;
  else
    g826 <= g13421;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g823 <= 0;
  else
    g823 <= gbuf71;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g853 <= 0;
  else
    g853 <= gbuf72;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g818 <= 0;
  else
    g818 <= g24300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g819 <= 0;
  else
    g819 <= g24301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g817 <= 0;
  else
    g817 <= g24302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g821 <= 0;
  else
    g821 <= g24303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g822 <= 0;
  else
    g822 <= g24304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g820 <= 0;
  else
    g820 <= g24305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g830 <= 0;
  else
    g830 <= g24306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g831 <= 0;
  else
    g831 <= g24307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g829 <= 0;
  else
    g829 <= g24308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g833 <= 0;
  else
    g833 <= g24309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g834 <= 0;
  else
    g834 <= g24310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g832 <= 0;
  else
    g832 <= g24311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g836 <= 0;
  else
    g836 <= g24312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g837 <= 0;
  else
    g837 <= g24313;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g835 <= 0;
  else
    g835 <= g24314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g839 <= 0;
  else
    g839 <= g24315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g840 <= 0;
  else
    g840 <= g24316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g838 <= 0;
  else
    g838 <= g24317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g842 <= 0;
  else
    g842 <= g24318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g843 <= 0;
  else
    g843 <= g24319;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g841 <= 0;
  else
    g841 <= g24320;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g845 <= 0;
  else
    g845 <= g24321;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g846 <= 0;
  else
    g846 <= g24322;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g844 <= 0;
  else
    g844 <= g24323;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g848 <= 0;
  else
    g848 <= g24324;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g849 <= 0;
  else
    g849 <= g24325;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g847 <= 0;
  else
    g847 <= g24326;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g851 <= 0;
  else
    g851 <= g24327;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g852 <= 0;
  else
    g852 <= g24328;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g850 <= 0;
  else
    g850 <= g24329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g857 <= 0;
  else
    g857 <= g26696;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g858 <= 0;
  else
    g858 <= g26697;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g856 <= 0;
  else
    g856 <= g26698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g860 <= 0;
  else
    g860 <= g26699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g861 <= 0;
  else
    g861 <= g26700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g859 <= 0;
  else
    g859 <= g26701;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g863 <= 0;
  else
    g863 <= g26702;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g864 <= 0;
  else
    g864 <= g26703;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g862 <= 0;
  else
    g862 <= g26704;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g866 <= 0;
  else
    g866 <= g26705;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g867 <= 0;
  else
    g867 <= g26706;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g865 <= 0;
  else
    g865 <= g26707;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g873 <= 0;
  else
    g873 <= g30521;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g876 <= 0;
  else
    g876 <= g30522;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g879 <= 0;
  else
    g879 <= g30523;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g918 <= 0;
  else
    g918 <= g30860;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g921 <= 0;
  else
    g921 <= g30861;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g924 <= 0;
  else
    g924 <= g30862;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g882 <= 0;
  else
    g882 <= g30854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g885 <= 0;
  else
    g885 <= g30855;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g888 <= 0;
  else
    g888 <= g30856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g927 <= 0;
  else
    g927 <= g30863;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g930 <= 0;
  else
    g930 <= g30864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g933 <= 0;
  else
    g933 <= g30865;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g891 <= 0;
  else
    g891 <= g30524;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g894 <= 0;
  else
    g894 <= g30525;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g897 <= 0;
  else
    g897 <= g30526;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g936 <= 0;
  else
    g936 <= g30530;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g939 <= 0;
  else
    g939 <= g30531;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g942 <= 0;
  else
    g942 <= g30532;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g900 <= 0;
  else
    g900 <= g30527;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g903 <= 0;
  else
    g903 <= g30528;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g906 <= 0;
  else
    g906 <= g30529;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g945 <= 0;
  else
    g945 <= g30533;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g948 <= 0;
  else
    g948 <= g30534;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g951 <= 0;
  else
    g951 <= g30535;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g909 <= 0;
  else
    g909 <= g30857;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g912 <= 0;
  else
    g912 <= g30858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g915 <= 0;
  else
    g915 <= g30859;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g954 <= 0;
  else
    g954 <= g30866;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g957 <= 0;
  else
    g957 <= g30867;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g960 <= 0;
  else
    g960 <= g30868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g780 <= 0;
  else
    g780 <= g25992;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g776 <= 0;
  else
    g776 <= g26695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g771 <= 0;
  else
    g771 <= g27198;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g767 <= 0;
  else
    g767 <= g27691;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g762 <= 0;
  else
    g762 <= g28232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g758 <= 0;
  else
    g758 <= g28678;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g753 <= 0;
  else
    g753 <= g29139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g749 <= 0;
  else
    g749 <= g29420;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g744 <= 0;
  else
    g744 <= g29634;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g740 <= 0;
  else
    g740 <= g29798;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g868 <= 0;
  else
    g868 <= g20559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g870 <= 0;
  else
    g870 <= gbuf73;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g869 <= 0;
  else
    g869 <= gbuf74;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g963 <= 0;
  else
    g963 <= g13422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1092 <= 0;
  else
    g1092 <= gbuf75;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1088 <= 0;
  else
    g1088 <= gbuf76;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g996 <= 0;
  else
    g996 <= g11523;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1041 <= 0;
  else
    g1041 <= g28233;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1030 <= 0;
  else
    g1030 <= g28234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1033 <= 0;
  else
    g1033 <= g28235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1056 <= 0;
  else
    g1056 <= g28236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1045 <= 0;
  else
    g1045 <= g28237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1048 <= 0;
  else
    g1048 <= g28238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1071 <= 0;
  else
    g1071 <= g28239;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1060 <= 0;
  else
    g1060 <= g28240;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1063 <= 0;
  else
    g1063 <= g28241;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1085 <= 0;
  else
    g1085 <= g28242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1075 <= 0;
  else
    g1075 <= g28243;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1078 <= 0;
  else
    g1078 <= g28244;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1095 <= 0;
  else
    g1095 <= g29421;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1098 <= 0;
  else
    g1098 <= g29422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1101 <= 0;
  else
    g1101 <= g29423;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1104 <= 0;
  else
    g1104 <= g29638;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1107 <= 0;
  else
    g1107 <= g29639;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1110 <= 0;
  else
    g1110 <= g29640;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1114 <= 0;
  else
    g1114 <= g29424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1115 <= 0;
  else
    g1115 <= g29425;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1113 <= 0;
  else
    g1113 <= g29426;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1116 <= 0;
  else
    g1116 <= g27692;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1119 <= 0;
  else
    g1119 <= g27693;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1122 <= 0;
  else
    g1122 <= g27694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1125 <= 0;
  else
    g1125 <= g27695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1128 <= 0;
  else
    g1128 <= g27696;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1131 <= 0;
  else
    g1131 <= g27697;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1135 <= 0;
  else
    g1135 <= g28679;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1136 <= 0;
  else
    g1136 <= g28680;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1134 <= 0;
  else
    g1134 <= g28681;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g999 <= 0;
  else
    g999 <= g29799;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1000 <= 0;
  else
    g1000 <= g29800;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1001 <= 0;
  else
    g1001 <= g29801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1002 <= 0;
  else
    g1002 <= g30869;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1003 <= 0;
  else
    g1003 <= g30870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1004 <= 0;
  else
    g1004 <= g30871;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1005 <= 0;
  else
    g1005 <= g30713;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1006 <= 0;
  else
    g1006 <= g30714;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1007 <= 0;
  else
    g1007 <= g30715;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1009 <= 0;
  else
    g1009 <= g29635;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1010 <= 0;
  else
    g1010 <= g29636;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1008 <= 0;
  else
    g1008 <= g29637;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1090 <= 0;
  else
    g1090 <= g27206;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1091 <= 0;
  else
    g1091 <= g27207;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1089 <= 0;
  else
    g1089 <= g27208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1137 <= 0;
  else
    g1137 <= g11536;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1138 <= 0;
  else
    g1138 <= gbuf77;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1139 <= 0;
  else
    g1139 <= g11537;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1140 <= 0;
  else
    g1140 <= gbuf78;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1141 <= 0;
  else
    g1141 <= g11538;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g966 <= 0;
  else
    g966 <= gbuf79;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g967 <= 0;
  else
    g967 <= g11518;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g968 <= 0;
  else
    g968 <= gbuf80;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g969 <= 0;
  else
    g969 <= g11519;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g970 <= 0;
  else
    g970 <= gbuf81;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g971 <= 0;
  else
    g971 <= g11520;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g972 <= 0;
  else
    g972 <= gbuf82;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g973 <= 0;
  else
    g973 <= g11521;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g974 <= 0;
  else
    g974 <= gbuf83;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g975 <= 0;
  else
    g975 <= g11522;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g976 <= 0;
  else
    g976 <= gbuf84;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g977 <= 0;
  else
    g977 <= g13423;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g978 <= 0;
  else
    g978 <= gbuf85;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g986 <= 0;
  else
    g986 <= g19024;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g992 <= 0;
  else
    g992 <= g27200;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g995 <= 0;
  else
    g995 <= g27201;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g984 <= 0;
  else
    g984 <= g27202;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g983 <= 0;
  else
    g983 <= g27203;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g982 <= 0;
  else
    g982 <= g27204;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g981 <= 0;
  else
    g981 <= g27205;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g991 <= 0;
  else
    g991 <= g19028;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g990 <= 0;
  else
    g990 <= g19027;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g989 <= 0;
  else
    g989 <= g19026;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g988 <= 0;
  else
    g988 <= g19025;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g987 <= 0;
  else
    g987 <= g25141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g985 <= 0;
  else
    g985 <= g27199;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1029 <= 0;
  else
    g1029 <= g11524;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1036 <= 0;
  else
    g1036 <= gbuf86;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1037 <= 0;
  else
    g1037 <= g11525;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1038 <= 0;
  else
    g1038 <= gbuf87;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1039 <= 0;
  else
    g1039 <= g11526;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1040 <= 0;
  else
    g1040 <= gbuf88;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1044 <= 0;
  else
    g1044 <= g11527;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1051 <= 0;
  else
    g1051 <= gbuf89;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1052 <= 0;
  else
    g1052 <= g11528;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1053 <= 0;
  else
    g1053 <= gbuf90;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1054 <= 0;
  else
    g1054 <= g11529;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1055 <= 0;
  else
    g1055 <= gbuf91;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1059 <= 0;
  else
    g1059 <= g11530;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1066 <= 0;
  else
    g1066 <= gbuf92;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1067 <= 0;
  else
    g1067 <= g11531;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1068 <= 0;
  else
    g1068 <= gbuf93;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1069 <= 0;
  else
    g1069 <= g11532;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1070 <= 0;
  else
    g1070 <= gbuf94;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1074 <= 0;
  else
    g1074 <= g11533;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1081 <= 0;
  else
    g1081 <= gbuf95;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1082 <= 0;
  else
    g1082 <= g11534;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1083 <= 0;
  else
    g1083 <= gbuf96;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1084 <= 0;
  else
    g1084 <= g11535;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1011 <= 0;
  else
    g1011 <= gbuf97;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1012 <= 0;
  else
    g1012 <= g13424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1018 <= 0;
  else
    g1018 <= gbuf98;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1024 <= 0;
  else
    g1024 <= gbuf99;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1231 <= 0;
  else
    g1231 <= g13435;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1237 <= 0;
  else
    g1237 <= gbuf100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1236 <= 0;
  else
    g1236 <= gbuf101;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1240 <= 0;
  else
    g1240 <= g23198;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1243 <= 0;
  else
    g1243 <= g20560;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1196 <= 0;
  else
    g1196 <= g20561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1199 <= 0;
  else
    g1199 <= g16469;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1209 <= 0;
  else
    g1209 <= gbuf102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1210 <= 0;
  else
    g1210 <= gbuf103;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1250 <= 0;
  else
    g1250 <= g11539;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1255 <= 0;
  else
    g1255 <= gbuf104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1256 <= 0;
  else
    g1256 <= g11542;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1257 <= 0;
  else
    g1257 <= gbuf105;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1258 <= 0;
  else
    g1258 <= g11543;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1259 <= 0;
  else
    g1259 <= gbuf106;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1260 <= 0;
  else
    g1260 <= g11544;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1251 <= 0;
  else
    g1251 <= gbuf107;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1252 <= 0;
  else
    g1252 <= g11540;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1253 <= 0;
  else
    g1253 <= gbuf108;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1254 <= 0;
  else
    g1254 <= g11541;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1176 <= 0;
  else
    g1176 <= gbuf109;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1161 <= 0;
  else
    g1161 <= g13425;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1168 <= 0;
  else
    g1168 <= gbuf110;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1172 <= 0;
  else
    g1172 <= gbuf111;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1173 <= 0;
  else
    g1173 <= g24333;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1174 <= 0;
  else
    g1174 <= g24334;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1175 <= 0;
  else
    g1175 <= g24335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1142 <= 0;
  else
    g1142 <= g25150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1145 <= 0;
  else
    g1145 <= g25142;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1148 <= 0;
  else
    g1148 <= g25143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1164 <= 0;
  else
    g1164 <= g25147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1165 <= 0;
  else
    g1165 <= g25148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1166 <= 0;
  else
    g1166 <= g25149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1167 <= 0;
  else
    g1167 <= g24330;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1171 <= 0;
  else
    g1171 <= g24331;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1151 <= 0;
  else
    g1151 <= g24332;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1152 <= 0;
  else
    g1152 <= g25144;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1155 <= 0;
  else
    g1155 <= g25145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1158 <= 0;
  else
    g1158 <= g25146;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1214 <= 0;
  else
    g1214 <= g16470;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1221 <= 0;
  else
    g1221 <= gbuf112;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1228 <= 0;
  else
    g1228 <= gbuf113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1229 <= 0;
  else
    g1229 <= g19033;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1230 <= 0;
  else
    g1230 <= gbuf114;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1234 <= 0;
  else
    g1234 <= g27217;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1235 <= 0;
  else
    g1235 <= g19034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1186 <= 0;
  else
    g1186 <= gbuf115;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1244 <= 0;
  else
    g1244 <= g19035;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1245 <= 0;
  else
    g1245 <= gbuf116;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1262 <= 0;
  else
    g1262 <= g28245;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1263 <= 0;
  else
    g1263 <= g28246;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1261 <= 0;
  else
    g1261 <= g28247;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1265 <= 0;
  else
    g1265 <= g28248;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1266 <= 0;
  else
    g1266 <= g28249;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1264 <= 0;
  else
    g1264 <= g28250;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1268 <= 0;
  else
    g1268 <= g28251;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1269 <= 0;
  else
    g1269 <= g28252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1267 <= 0;
  else
    g1267 <= g28253;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1271 <= 0;
  else
    g1271 <= g28254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1272 <= 0;
  else
    g1272 <= g28255;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1270 <= 0;
  else
    g1270 <= g28256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1273 <= 0;
  else
    g1273 <= g25994;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1276 <= 0;
  else
    g1276 <= g25995;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1279 <= 0;
  else
    g1279 <= g25996;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1282 <= 0;
  else
    g1282 <= g25997;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1285 <= 0;
  else
    g1285 <= g25998;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1288 <= 0;
  else
    g1288 <= g25999;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1300 <= 0;
  else
    g1300 <= g29143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1303 <= 0;
  else
    g1303 <= g29144;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1306 <= 0;
  else
    g1306 <= g29145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1291 <= 0;
  else
    g1291 <= g29140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1294 <= 0;
  else
    g1294 <= g29141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1297 <= 0;
  else
    g1297 <= g29142;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1177 <= 0;
  else
    g1177 <= g27209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1180 <= 0;
  else
    g1180 <= g27210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1183 <= 0;
  else
    g1183 <= g27211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1192 <= 0;
  else
    g1192 <= g8293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1193 <= 0;
  else
    g1193 <= g24336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1194 <= 0;
  else
    g1194 <= g19029;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1195 <= 0;
  else
    g1195 <= g19030;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1200 <= 0;
  else
    g1200 <= g19031;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1201 <= 0;
  else
    g1201 <= g19032;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1202 <= 0;
  else
    g1202 <= g27216;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1203 <= 0;
  else
    g1203 <= g27215;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1204 <= 0;
  else
    g1204 <= g27214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1205 <= 0;
  else
    g1205 <= g27213;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1206 <= 0;
  else
    g1206 <= g27212;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1211 <= 0;
  else
    g1211 <= gbuf117;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1215 <= 0;
  else
    g1215 <= g13426;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1216 <= 0;
  else
    g1216 <= g13427;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1217 <= 0;
  else
    g1217 <= g13428;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1218 <= 0;
  else
    g1218 <= g13429;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1219 <= 0;
  else
    g1219 <= g13430;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1220 <= 0;
  else
    g1220 <= g13431;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1222 <= 0;
  else
    g1222 <= g13432;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1223 <= 0;
  else
    g1223 <= g13433;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1224 <= 0;
  else
    g1224 <= g25993;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1227 <= 0;
  else
    g1227 <= g13434;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1309 <= 0;
  else
    g1309 <= g13436;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1312 <= 0;
  else
    g1312 <= gbuf118;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1315 <= 0;
  else
    g1315 <= gbuf119;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1316 <= 0;
  else
    g1316 <= g20562;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1345 <= 0;
  else
    g1345 <= g21944;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1326 <= 0;
  else
    g1326 <= g23199;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1319 <= 0;
  else
    g1319 <= g24337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1339 <= 0;
  else
    g1339 <= g25151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1332 <= 0;
  else
    g1332 <= g26000;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1346 <= 0;
  else
    g1346 <= g26708;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1358 <= 0;
  else
    g1358 <= g27218;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1352 <= 0;
  else
    g1352 <= g27698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1365 <= 0;
  else
    g1365 <= g28257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1372 <= 0;
  else
    g1372 <= g28682;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1378 <= 0;
  else
    g1378 <= g29146;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1385 <= 0;
  else
    g1385 <= g23200;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1386 <= 0;
  else
    g1386 <= g23201;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1384 <= 0;
  else
    g1384 <= g23202;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1388 <= 0;
  else
    g1388 <= g23203;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1389 <= 0;
  else
    g1389 <= g23204;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1387 <= 0;
  else
    g1387 <= g23205;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1391 <= 0;
  else
    g1391 <= g23206;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1392 <= 0;
  else
    g1392 <= g23207;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1390 <= 0;
  else
    g1390 <= g23208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1394 <= 0;
  else
    g1394 <= g23209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1395 <= 0;
  else
    g1395 <= g23210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1393 <= 0;
  else
    g1393 <= g23211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1397 <= 0;
  else
    g1397 <= g23212;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1398 <= 0;
  else
    g1398 <= g23213;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1396 <= 0;
  else
    g1396 <= g23214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1400 <= 0;
  else
    g1400 <= g23215;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1401 <= 0;
  else
    g1401 <= g23216;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1399 <= 0;
  else
    g1399 <= g23217;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1403 <= 0;
  else
    g1403 <= g23218;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1404 <= 0;
  else
    g1404 <= g23219;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1402 <= 0;
  else
    g1402 <= g23220;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1406 <= 0;
  else
    g1406 <= g23221;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1407 <= 0;
  else
    g1407 <= g23222;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1405 <= 0;
  else
    g1405 <= g23223;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1409 <= 0;
  else
    g1409 <= g23224;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1410 <= 0;
  else
    g1410 <= g23225;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1408 <= 0;
  else
    g1408 <= g23226;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1412 <= 0;
  else
    g1412 <= g23227;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1413 <= 0;
  else
    g1413 <= g23228;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1411 <= 0;
  else
    g1411 <= g23229;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1415 <= 0;
  else
    g1415 <= g23230;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1416 <= 0;
  else
    g1416 <= g23231;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1414 <= 0;
  else
    g1414 <= g23232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1418 <= 0;
  else
    g1418 <= g23233;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1419 <= 0;
  else
    g1419 <= g23234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1417 <= 0;
  else
    g1417 <= g23235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1421 <= 0;
  else
    g1421 <= g26709;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1422 <= 0;
  else
    g1422 <= g26710;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1420 <= 0;
  else
    g1420 <= g26711;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1424 <= 0;
  else
    g1424 <= g24338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1425 <= 0;
  else
    g1425 <= g24339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1423 <= 0;
  else
    g1423 <= g24340;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1520 <= 0;
  else
    g1520 <= g13437;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1517 <= 0;
  else
    g1517 <= gbuf120;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1547 <= 0;
  else
    g1547 <= gbuf121;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1512 <= 0;
  else
    g1512 <= g24341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1513 <= 0;
  else
    g1513 <= g24342;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1511 <= 0;
  else
    g1511 <= g24343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1515 <= 0;
  else
    g1515 <= g24344;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1516 <= 0;
  else
    g1516 <= g24345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1514 <= 0;
  else
    g1514 <= g24346;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1524 <= 0;
  else
    g1524 <= g24347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1525 <= 0;
  else
    g1525 <= g24348;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1523 <= 0;
  else
    g1523 <= g24349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1527 <= 0;
  else
    g1527 <= g24350;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1528 <= 0;
  else
    g1528 <= g24351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1526 <= 0;
  else
    g1526 <= g24352;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1530 <= 0;
  else
    g1530 <= g24353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1531 <= 0;
  else
    g1531 <= g24354;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1529 <= 0;
  else
    g1529 <= g24355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1533 <= 0;
  else
    g1533 <= g24356;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1534 <= 0;
  else
    g1534 <= g24357;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1532 <= 0;
  else
    g1532 <= g24358;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1536 <= 0;
  else
    g1536 <= g24359;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1537 <= 0;
  else
    g1537 <= g24360;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1535 <= 0;
  else
    g1535 <= g24361;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1539 <= 0;
  else
    g1539 <= g24362;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1540 <= 0;
  else
    g1540 <= g24363;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1538 <= 0;
  else
    g1538 <= g24364;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1542 <= 0;
  else
    g1542 <= g24365;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1543 <= 0;
  else
    g1543 <= g24366;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1541 <= 0;
  else
    g1541 <= g24367;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1545 <= 0;
  else
    g1545 <= g24368;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1546 <= 0;
  else
    g1546 <= g24369;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1544 <= 0;
  else
    g1544 <= g24370;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1551 <= 0;
  else
    g1551 <= g26713;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1552 <= 0;
  else
    g1552 <= g26714;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1550 <= 0;
  else
    g1550 <= g26715;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1554 <= 0;
  else
    g1554 <= g26716;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1555 <= 0;
  else
    g1555 <= g26717;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1553 <= 0;
  else
    g1553 <= g26718;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1557 <= 0;
  else
    g1557 <= g26719;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1558 <= 0;
  else
    g1558 <= g26720;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1556 <= 0;
  else
    g1556 <= g26721;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1560 <= 0;
  else
    g1560 <= g26722;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1561 <= 0;
  else
    g1561 <= g26723;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1559 <= 0;
  else
    g1559 <= g26724;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1567 <= 0;
  else
    g1567 <= g30536;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1570 <= 0;
  else
    g1570 <= g30537;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1573 <= 0;
  else
    g1573 <= g30538;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1612 <= 0;
  else
    g1612 <= g30878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1615 <= 0;
  else
    g1615 <= g30879;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1618 <= 0;
  else
    g1618 <= g30880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1576 <= 0;
  else
    g1576 <= g30872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1579 <= 0;
  else
    g1579 <= g30873;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1582 <= 0;
  else
    g1582 <= g30874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1621 <= 0;
  else
    g1621 <= g30881;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1624 <= 0;
  else
    g1624 <= g30882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1627 <= 0;
  else
    g1627 <= g30883;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1585 <= 0;
  else
    g1585 <= g30539;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1588 <= 0;
  else
    g1588 <= g30540;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1591 <= 0;
  else
    g1591 <= g30541;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1630 <= 0;
  else
    g1630 <= g30545;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1633 <= 0;
  else
    g1633 <= g30546;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1636 <= 0;
  else
    g1636 <= g30547;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1594 <= 0;
  else
    g1594 <= g30542;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1597 <= 0;
  else
    g1597 <= g30543;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1600 <= 0;
  else
    g1600 <= g30544;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1639 <= 0;
  else
    g1639 <= g30548;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1642 <= 0;
  else
    g1642 <= g30549;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1645 <= 0;
  else
    g1645 <= g30550;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1603 <= 0;
  else
    g1603 <= g30875;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1606 <= 0;
  else
    g1606 <= g30876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1609 <= 0;
  else
    g1609 <= g30877;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1648 <= 0;
  else
    g1648 <= g30884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1651 <= 0;
  else
    g1651 <= g30885;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1654 <= 0;
  else
    g1654 <= g30886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1466 <= 0;
  else
    g1466 <= g26001;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1462 <= 0;
  else
    g1462 <= g26712;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1457 <= 0;
  else
    g1457 <= g27219;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1453 <= 0;
  else
    g1453 <= g27699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1448 <= 0;
  else
    g1448 <= g28258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1444 <= 0;
  else
    g1444 <= g28683;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1439 <= 0;
  else
    g1439 <= g29147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1435 <= 0;
  else
    g1435 <= g29427;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1430 <= 0;
  else
    g1430 <= g29641;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1426 <= 0;
  else
    g1426 <= g29802;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1562 <= 0;
  else
    g1562 <= g20563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1564 <= 0;
  else
    g1564 <= gbuf122;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1563 <= 0;
  else
    g1563 <= gbuf123;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1657 <= 0;
  else
    g1657 <= g13438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1786 <= 0;
  else
    g1786 <= gbuf124;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1782 <= 0;
  else
    g1782 <= gbuf125;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1690 <= 0;
  else
    g1690 <= g11550;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1735 <= 0;
  else
    g1735 <= g28259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1724 <= 0;
  else
    g1724 <= g28260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1727 <= 0;
  else
    g1727 <= g28261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1750 <= 0;
  else
    g1750 <= g28262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1739 <= 0;
  else
    g1739 <= g28263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1742 <= 0;
  else
    g1742 <= g28264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1765 <= 0;
  else
    g1765 <= g28265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1754 <= 0;
  else
    g1754 <= g28266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1757 <= 0;
  else
    g1757 <= g28267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1779 <= 0;
  else
    g1779 <= g28268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1769 <= 0;
  else
    g1769 <= g28269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1772 <= 0;
  else
    g1772 <= g28270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1789 <= 0;
  else
    g1789 <= g29434;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1792 <= 0;
  else
    g1792 <= g29435;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1795 <= 0;
  else
    g1795 <= g29436;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1798 <= 0;
  else
    g1798 <= g29645;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1801 <= 0;
  else
    g1801 <= g29646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1804 <= 0;
  else
    g1804 <= g29647;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1808 <= 0;
  else
    g1808 <= g29437;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1809 <= 0;
  else
    g1809 <= g29438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1807 <= 0;
  else
    g1807 <= g29439;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1810 <= 0;
  else
    g1810 <= g27700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1813 <= 0;
  else
    g1813 <= g27701;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1816 <= 0;
  else
    g1816 <= g27702;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1819 <= 0;
  else
    g1819 <= g27703;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1822 <= 0;
  else
    g1822 <= g27704;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1825 <= 0;
  else
    g1825 <= g27705;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1829 <= 0;
  else
    g1829 <= g28684;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1830 <= 0;
  else
    g1830 <= g28685;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1828 <= 0;
  else
    g1828 <= g28686;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1693 <= 0;
  else
    g1693 <= g29803;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1694 <= 0;
  else
    g1694 <= g29804;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1695 <= 0;
  else
    g1695 <= g29805;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1696 <= 0;
  else
    g1696 <= g30887;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1697 <= 0;
  else
    g1697 <= g30888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1698 <= 0;
  else
    g1698 <= g30889;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1699 <= 0;
  else
    g1699 <= g30716;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1700 <= 0;
  else
    g1700 <= g30717;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1701 <= 0;
  else
    g1701 <= g30718;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1703 <= 0;
  else
    g1703 <= g29642;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1704 <= 0;
  else
    g1704 <= g29643;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1702 <= 0;
  else
    g1702 <= g29644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1784 <= 0;
  else
    g1784 <= g27221;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1785 <= 0;
  else
    g1785 <= g27222;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1783 <= 0;
  else
    g1783 <= g27223;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1831 <= 0;
  else
    g1831 <= g11563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1832 <= 0;
  else
    g1832 <= gbuf126;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1833 <= 0;
  else
    g1833 <= g11564;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1834 <= 0;
  else
    g1834 <= gbuf127;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1835 <= 0;
  else
    g1835 <= g11565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1660 <= 0;
  else
    g1660 <= gbuf128;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1661 <= 0;
  else
    g1661 <= g11545;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1662 <= 0;
  else
    g1662 <= gbuf129;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1663 <= 0;
  else
    g1663 <= g11546;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1664 <= 0;
  else
    g1664 <= gbuf130;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1665 <= 0;
  else
    g1665 <= g11547;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1666 <= 0;
  else
    g1666 <= gbuf131;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1667 <= 0;
  else
    g1667 <= g11548;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1668 <= 0;
  else
    g1668 <= gbuf132;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1669 <= 0;
  else
    g1669 <= g11549;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1670 <= 0;
  else
    g1670 <= gbuf133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1671 <= 0;
  else
    g1671 <= g13439;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1672 <= 0;
  else
    g1672 <= gbuf134;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1680 <= 0;
  else
    g1680 <= g19036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1686 <= 0;
  else
    g1686 <= g29428;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1689 <= 0;
  else
    g1689 <= g29429;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1678 <= 0;
  else
    g1678 <= g29430;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1677 <= 0;
  else
    g1677 <= g29431;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1676 <= 0;
  else
    g1676 <= g29432;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1675 <= 0;
  else
    g1675 <= g29433;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1685 <= 0;
  else
    g1685 <= g19040;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1684 <= 0;
  else
    g1684 <= g19039;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1683 <= 0;
  else
    g1683 <= g19038;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1682 <= 0;
  else
    g1682 <= g19037;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1681 <= 0;
  else
    g1681 <= g25152;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1679 <= 0;
  else
    g1679 <= g27220;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1723 <= 0;
  else
    g1723 <= g11551;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1730 <= 0;
  else
    g1730 <= gbuf135;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1731 <= 0;
  else
    g1731 <= g11552;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1732 <= 0;
  else
    g1732 <= gbuf136;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1733 <= 0;
  else
    g1733 <= g11553;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1734 <= 0;
  else
    g1734 <= gbuf137;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1738 <= 0;
  else
    g1738 <= g11554;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1745 <= 0;
  else
    g1745 <= gbuf138;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1746 <= 0;
  else
    g1746 <= g11555;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1747 <= 0;
  else
    g1747 <= gbuf139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1748 <= 0;
  else
    g1748 <= g11556;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1749 <= 0;
  else
    g1749 <= gbuf140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1753 <= 0;
  else
    g1753 <= g11557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1760 <= 0;
  else
    g1760 <= gbuf141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1761 <= 0;
  else
    g1761 <= g11558;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1762 <= 0;
  else
    g1762 <= gbuf142;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1763 <= 0;
  else
    g1763 <= g11559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1764 <= 0;
  else
    g1764 <= gbuf143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1768 <= 0;
  else
    g1768 <= g11560;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1775 <= 0;
  else
    g1775 <= gbuf144;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1776 <= 0;
  else
    g1776 <= g11561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1777 <= 0;
  else
    g1777 <= gbuf145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1778 <= 0;
  else
    g1778 <= g11562;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1705 <= 0;
  else
    g1705 <= gbuf146;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1706 <= 0;
  else
    g1706 <= g13440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1712 <= 0;
  else
    g1712 <= gbuf147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1718 <= 0;
  else
    g1718 <= gbuf148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1925 <= 0;
  else
    g1925 <= g13451;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1931 <= 0;
  else
    g1931 <= gbuf149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1930 <= 0;
  else
    g1930 <= gbuf150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1934 <= 0;
  else
    g1934 <= g23236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1937 <= 0;
  else
    g1937 <= g20564;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1890 <= 0;
  else
    g1890 <= g20565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1893 <= 0;
  else
    g1893 <= g16471;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1903 <= 0;
  else
    g1903 <= gbuf151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1904 <= 0;
  else
    g1904 <= gbuf152;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1944 <= 0;
  else
    g1944 <= g11566;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1949 <= 0;
  else
    g1949 <= gbuf153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1950 <= 0;
  else
    g1950 <= g11569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1951 <= 0;
  else
    g1951 <= gbuf154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1952 <= 0;
  else
    g1952 <= g11570;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1953 <= 0;
  else
    g1953 <= gbuf155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1954 <= 0;
  else
    g1954 <= g11571;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1945 <= 0;
  else
    g1945 <= gbuf156;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1946 <= 0;
  else
    g1946 <= g11567;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1947 <= 0;
  else
    g1947 <= gbuf157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1948 <= 0;
  else
    g1948 <= g11568;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1870 <= 0;
  else
    g1870 <= gbuf158;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1855 <= 0;
  else
    g1855 <= g13441;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1862 <= 0;
  else
    g1862 <= gbuf159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1866 <= 0;
  else
    g1866 <= gbuf160;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1867 <= 0;
  else
    g1867 <= g24374;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1868 <= 0;
  else
    g1868 <= g24375;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1869 <= 0;
  else
    g1869 <= g24376;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1836 <= 0;
  else
    g1836 <= g25161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1839 <= 0;
  else
    g1839 <= g25153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1842 <= 0;
  else
    g1842 <= g25154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1858 <= 0;
  else
    g1858 <= g25158;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1859 <= 0;
  else
    g1859 <= g25159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1860 <= 0;
  else
    g1860 <= g25160;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1861 <= 0;
  else
    g1861 <= g24371;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1865 <= 0;
  else
    g1865 <= g24372;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1845 <= 0;
  else
    g1845 <= g24373;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1846 <= 0;
  else
    g1846 <= g25155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1849 <= 0;
  else
    g1849 <= g25156;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1852 <= 0;
  else
    g1852 <= g25157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1908 <= 0;
  else
    g1908 <= g16472;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1915 <= 0;
  else
    g1915 <= gbuf161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1922 <= 0;
  else
    g1922 <= gbuf162;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1923 <= 0;
  else
    g1923 <= g19045;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1924 <= 0;
  else
    g1924 <= gbuf163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1928 <= 0;
  else
    g1928 <= g29445;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1929 <= 0;
  else
    g1929 <= g19046;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1880 <= 0;
  else
    g1880 <= gbuf164;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1938 <= 0;
  else
    g1938 <= g19047;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1939 <= 0;
  else
    g1939 <= gbuf165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1956 <= 0;
  else
    g1956 <= g28271;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1957 <= 0;
  else
    g1957 <= g28272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1955 <= 0;
  else
    g1955 <= g28273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1959 <= 0;
  else
    g1959 <= g28274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1960 <= 0;
  else
    g1960 <= g28275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1958 <= 0;
  else
    g1958 <= g28276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1962 <= 0;
  else
    g1962 <= g28277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1963 <= 0;
  else
    g1963 <= g28278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1961 <= 0;
  else
    g1961 <= g28279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1965 <= 0;
  else
    g1965 <= g28280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1966 <= 0;
  else
    g1966 <= g28281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1964 <= 0;
  else
    g1964 <= g28282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1967 <= 0;
  else
    g1967 <= g26003;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1970 <= 0;
  else
    g1970 <= g26004;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1973 <= 0;
  else
    g1973 <= g26005;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1976 <= 0;
  else
    g1976 <= g26006;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1979 <= 0;
  else
    g1979 <= g26007;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1982 <= 0;
  else
    g1982 <= g26008;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1994 <= 0;
  else
    g1994 <= g29151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1997 <= 0;
  else
    g1997 <= g29152;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2000 <= 0;
  else
    g2000 <= g29153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1985 <= 0;
  else
    g1985 <= g29148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1988 <= 0;
  else
    g1988 <= g29149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1991 <= 0;
  else
    g1991 <= g29150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1871 <= 0;
  else
    g1871 <= g27224;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1874 <= 0;
  else
    g1874 <= g27225;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1877 <= 0;
  else
    g1877 <= g27226;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1886 <= 0;
  else
    g1886 <= g8302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1887 <= 0;
  else
    g1887 <= g24377;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1888 <= 0;
  else
    g1888 <= g19041;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1889 <= 0;
  else
    g1889 <= g19042;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1894 <= 0;
  else
    g1894 <= g19043;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1895 <= 0;
  else
    g1895 <= g19044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1896 <= 0;
  else
    g1896 <= g29444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1897 <= 0;
  else
    g1897 <= g29443;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1898 <= 0;
  else
    g1898 <= g29442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1899 <= 0;
  else
    g1899 <= g29441;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1900 <= 0;
  else
    g1900 <= g29440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1905 <= 0;
  else
    g1905 <= gbuf166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1909 <= 0;
  else
    g1909 <= g13442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1910 <= 0;
  else
    g1910 <= g13443;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1911 <= 0;
  else
    g1911 <= g13444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1912 <= 0;
  else
    g1912 <= g13445;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1913 <= 0;
  else
    g1913 <= g13446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1914 <= 0;
  else
    g1914 <= g13447;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1916 <= 0;
  else
    g1916 <= g13448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1917 <= 0;
  else
    g1917 <= g13449;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1918 <= 0;
  else
    g1918 <= g26002;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1921 <= 0;
  else
    g1921 <= g13450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2003 <= 0;
  else
    g2003 <= g13452;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2006 <= 0;
  else
    g2006 <= gbuf167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2009 <= 0;
  else
    g2009 <= gbuf168;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2010 <= 0;
  else
    g2010 <= g20566;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2039 <= 0;
  else
    g2039 <= g21945;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2020 <= 0;
  else
    g2020 <= g23237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2013 <= 0;
  else
    g2013 <= g24378;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2033 <= 0;
  else
    g2033 <= g25162;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2026 <= 0;
  else
    g2026 <= g26009;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2040 <= 0;
  else
    g2040 <= g26725;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2052 <= 0;
  else
    g2052 <= g27227;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2046 <= 0;
  else
    g2046 <= g27706;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2059 <= 0;
  else
    g2059 <= g28283;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2066 <= 0;
  else
    g2066 <= g28687;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2072 <= 0;
  else
    g2072 <= g29154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2079 <= 0;
  else
    g2079 <= g23238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2080 <= 0;
  else
    g2080 <= g23239;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2078 <= 0;
  else
    g2078 <= g23240;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2082 <= 0;
  else
    g2082 <= g23241;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2083 <= 0;
  else
    g2083 <= g23242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2081 <= 0;
  else
    g2081 <= g23243;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2085 <= 0;
  else
    g2085 <= g23244;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2086 <= 0;
  else
    g2086 <= g23245;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2084 <= 0;
  else
    g2084 <= g23246;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2088 <= 0;
  else
    g2088 <= g23247;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2089 <= 0;
  else
    g2089 <= g23248;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2087 <= 0;
  else
    g2087 <= g23249;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2091 <= 0;
  else
    g2091 <= g23250;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2092 <= 0;
  else
    g2092 <= g23251;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2090 <= 0;
  else
    g2090 <= g23252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2094 <= 0;
  else
    g2094 <= g23253;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2095 <= 0;
  else
    g2095 <= g23254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2093 <= 0;
  else
    g2093 <= g23255;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2097 <= 0;
  else
    g2097 <= g23256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2098 <= 0;
  else
    g2098 <= g23257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2096 <= 0;
  else
    g2096 <= g23258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2100 <= 0;
  else
    g2100 <= g23259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2101 <= 0;
  else
    g2101 <= g23260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2099 <= 0;
  else
    g2099 <= g23261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2103 <= 0;
  else
    g2103 <= g23262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2104 <= 0;
  else
    g2104 <= g23263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2102 <= 0;
  else
    g2102 <= g23264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2106 <= 0;
  else
    g2106 <= g23265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2107 <= 0;
  else
    g2107 <= g23266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2105 <= 0;
  else
    g2105 <= g23267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2109 <= 0;
  else
    g2109 <= g23268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2110 <= 0;
  else
    g2110 <= g23269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2108 <= 0;
  else
    g2108 <= g23270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2112 <= 0;
  else
    g2112 <= g23271;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2113 <= 0;
  else
    g2113 <= g23272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2111 <= 0;
  else
    g2111 <= g23273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2115 <= 0;
  else
    g2115 <= g26726;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2116 <= 0;
  else
    g2116 <= g26727;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2114 <= 0;
  else
    g2114 <= g26728;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2118 <= 0;
  else
    g2118 <= g24379;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2119 <= 0;
  else
    g2119 <= g24380;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2117 <= 0;
  else
    g2117 <= g24381;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2214 <= 0;
  else
    g2214 <= g13453;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2211 <= 0;
  else
    g2211 <= gbuf169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2241 <= 0;
  else
    g2241 <= gbuf170;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2206 <= 0;
  else
    g2206 <= g24382;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2207 <= 0;
  else
    g2207 <= g24383;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2205 <= 0;
  else
    g2205 <= g24384;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2209 <= 0;
  else
    g2209 <= g24385;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2210 <= 0;
  else
    g2210 <= g24386;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2208 <= 0;
  else
    g2208 <= g24387;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2218 <= 0;
  else
    g2218 <= g24388;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2219 <= 0;
  else
    g2219 <= g24389;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2217 <= 0;
  else
    g2217 <= g24390;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2221 <= 0;
  else
    g2221 <= g24391;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2222 <= 0;
  else
    g2222 <= g24392;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2220 <= 0;
  else
    g2220 <= g24393;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2224 <= 0;
  else
    g2224 <= g24394;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2225 <= 0;
  else
    g2225 <= g24395;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2223 <= 0;
  else
    g2223 <= g24396;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2227 <= 0;
  else
    g2227 <= g24397;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2228 <= 0;
  else
    g2228 <= g24398;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2226 <= 0;
  else
    g2226 <= g24399;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2230 <= 0;
  else
    g2230 <= g24400;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2231 <= 0;
  else
    g2231 <= g24401;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2229 <= 0;
  else
    g2229 <= g24402;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2233 <= 0;
  else
    g2233 <= g24403;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2234 <= 0;
  else
    g2234 <= g24404;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2232 <= 0;
  else
    g2232 <= g24405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2236 <= 0;
  else
    g2236 <= g24406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2237 <= 0;
  else
    g2237 <= g24407;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2235 <= 0;
  else
    g2235 <= g24408;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2239 <= 0;
  else
    g2239 <= g24409;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2240 <= 0;
  else
    g2240 <= g24410;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2238 <= 0;
  else
    g2238 <= g24411;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2245 <= 0;
  else
    g2245 <= g26730;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2246 <= 0;
  else
    g2246 <= g26731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2244 <= 0;
  else
    g2244 <= g26732;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2248 <= 0;
  else
    g2248 <= g26733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2249 <= 0;
  else
    g2249 <= g26734;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2247 <= 0;
  else
    g2247 <= g26735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2251 <= 0;
  else
    g2251 <= g26736;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2252 <= 0;
  else
    g2252 <= g26737;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2250 <= 0;
  else
    g2250 <= g26738;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2254 <= 0;
  else
    g2254 <= g26739;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2255 <= 0;
  else
    g2255 <= g26740;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2253 <= 0;
  else
    g2253 <= g26741;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2261 <= 0;
  else
    g2261 <= g30551;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2264 <= 0;
  else
    g2264 <= g30552;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2267 <= 0;
  else
    g2267 <= g30553;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2306 <= 0;
  else
    g2306 <= g30896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2309 <= 0;
  else
    g2309 <= g30897;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2312 <= 0;
  else
    g2312 <= g30898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2270 <= 0;
  else
    g2270 <= g30890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2273 <= 0;
  else
    g2273 <= g30891;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2276 <= 0;
  else
    g2276 <= g30892;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2315 <= 0;
  else
    g2315 <= g30899;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2318 <= 0;
  else
    g2318 <= g30900;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2321 <= 0;
  else
    g2321 <= g30901;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2279 <= 0;
  else
    g2279 <= g30554;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2282 <= 0;
  else
    g2282 <= g30555;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2285 <= 0;
  else
    g2285 <= g30556;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2324 <= 0;
  else
    g2324 <= g30560;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2327 <= 0;
  else
    g2327 <= g30561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2330 <= 0;
  else
    g2330 <= g30562;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2288 <= 0;
  else
    g2288 <= g30557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2291 <= 0;
  else
    g2291 <= g30558;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2294 <= 0;
  else
    g2294 <= g30559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2333 <= 0;
  else
    g2333 <= g30563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2336 <= 0;
  else
    g2336 <= g30564;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2339 <= 0;
  else
    g2339 <= g30565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2297 <= 0;
  else
    g2297 <= g30893;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2300 <= 0;
  else
    g2300 <= g30894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2303 <= 0;
  else
    g2303 <= g30895;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2342 <= 0;
  else
    g2342 <= g30902;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2345 <= 0;
  else
    g2345 <= g30903;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2348 <= 0;
  else
    g2348 <= g30904;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2160 <= 0;
  else
    g2160 <= g26010;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2156 <= 0;
  else
    g2156 <= g26729;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2151 <= 0;
  else
    g2151 <= g27228;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2147 <= 0;
  else
    g2147 <= g27707;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2142 <= 0;
  else
    g2142 <= g28284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2138 <= 0;
  else
    g2138 <= g28688;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2133 <= 0;
  else
    g2133 <= g29155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2129 <= 0;
  else
    g2129 <= g29446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2124 <= 0;
  else
    g2124 <= g29648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2120 <= 0;
  else
    g2120 <= g29806;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2256 <= 0;
  else
    g2256 <= g20567;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2258 <= 0;
  else
    g2258 <= gbuf171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2257 <= 0;
  else
    g2257 <= gbuf172;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2351 <= 0;
  else
    g2351 <= g13454;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2480 <= 0;
  else
    g2480 <= gbuf173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2476 <= 0;
  else
    g2476 <= gbuf174;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2384 <= 0;
  else
    g2384 <= g11577;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2429 <= 0;
  else
    g2429 <= g28285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2418 <= 0;
  else
    g2418 <= g28286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2421 <= 0;
  else
    g2421 <= g28287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2444 <= 0;
  else
    g2444 <= g28288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2433 <= 0;
  else
    g2433 <= g28289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2436 <= 0;
  else
    g2436 <= g28290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2459 <= 0;
  else
    g2459 <= g28291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2448 <= 0;
  else
    g2448 <= g28292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2451 <= 0;
  else
    g2451 <= g28293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2473 <= 0;
  else
    g2473 <= g28294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2463 <= 0;
  else
    g2463 <= g28295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2466 <= 0;
  else
    g2466 <= g28296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2483 <= 0;
  else
    g2483 <= g29447;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2486 <= 0;
  else
    g2486 <= g29448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2489 <= 0;
  else
    g2489 <= g29449;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2492 <= 0;
  else
    g2492 <= g29652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2495 <= 0;
  else
    g2495 <= g29653;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2498 <= 0;
  else
    g2498 <= g29654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2502 <= 0;
  else
    g2502 <= g29450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2503 <= 0;
  else
    g2503 <= g29451;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2501 <= 0;
  else
    g2501 <= g29452;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2504 <= 0;
  else
    g2504 <= g27708;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2507 <= 0;
  else
    g2507 <= g27709;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2510 <= 0;
  else
    g2510 <= g27710;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2513 <= 0;
  else
    g2513 <= g27711;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2516 <= 0;
  else
    g2516 <= g27712;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2519 <= 0;
  else
    g2519 <= g27713;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2523 <= 0;
  else
    g2523 <= g28689;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2524 <= 0;
  else
    g2524 <= g28690;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2522 <= 0;
  else
    g2522 <= g28691;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2387 <= 0;
  else
    g2387 <= g29807;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2388 <= 0;
  else
    g2388 <= g29808;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2389 <= 0;
  else
    g2389 <= g29809;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2390 <= 0;
  else
    g2390 <= g30905;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2391 <= 0;
  else
    g2391 <= g30906;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2392 <= 0;
  else
    g2392 <= g30907;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2393 <= 0;
  else
    g2393 <= g30719;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2394 <= 0;
  else
    g2394 <= g30720;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2395 <= 0;
  else
    g2395 <= g30721;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2397 <= 0;
  else
    g2397 <= g29649;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2398 <= 0;
  else
    g2398 <= g29650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2396 <= 0;
  else
    g2396 <= g29651;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2478 <= 0;
  else
    g2478 <= g27230;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2479 <= 0;
  else
    g2479 <= g27231;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2477 <= 0;
  else
    g2477 <= g27232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2525 <= 0;
  else
    g2525 <= g11590;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2526 <= 0;
  else
    g2526 <= gbuf175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2527 <= 0;
  else
    g2527 <= g11591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2528 <= 0;
  else
    g2528 <= gbuf176;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2529 <= 0;
  else
    g2529 <= g11592;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2354 <= 0;
  else
    g2354 <= gbuf177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2355 <= 0;
  else
    g2355 <= g11572;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2356 <= 0;
  else
    g2356 <= gbuf178;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2357 <= 0;
  else
    g2357 <= g11573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2358 <= 0;
  else
    g2358 <= gbuf179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2359 <= 0;
  else
    g2359 <= g11574;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2360 <= 0;
  else
    g2360 <= gbuf180;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2361 <= 0;
  else
    g2361 <= g11575;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2362 <= 0;
  else
    g2362 <= gbuf181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2363 <= 0;
  else
    g2363 <= g11576;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2364 <= 0;
  else
    g2364 <= gbuf182;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2365 <= 0;
  else
    g2365 <= g13455;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2366 <= 0;
  else
    g2366 <= gbuf183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2374 <= 0;
  else
    g2374 <= g19048;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2380 <= 0;
  else
    g2380 <= g30314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2383 <= 0;
  else
    g2383 <= g30315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2372 <= 0;
  else
    g2372 <= g30316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2371 <= 0;
  else
    g2371 <= g30317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2370 <= 0;
  else
    g2370 <= g30318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2369 <= 0;
  else
    g2369 <= g30319;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2379 <= 0;
  else
    g2379 <= g19052;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2378 <= 0;
  else
    g2378 <= g19051;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2377 <= 0;
  else
    g2377 <= g19050;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2376 <= 0;
  else
    g2376 <= g19049;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2375 <= 0;
  else
    g2375 <= g25163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2373 <= 0;
  else
    g2373 <= g27229;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2417 <= 0;
  else
    g2417 <= g11578;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2424 <= 0;
  else
    g2424 <= gbuf184;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2425 <= 0;
  else
    g2425 <= g11579;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2426 <= 0;
  else
    g2426 <= gbuf185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2427 <= 0;
  else
    g2427 <= g11580;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2428 <= 0;
  else
    g2428 <= gbuf186;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2432 <= 0;
  else
    g2432 <= g11581;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2439 <= 0;
  else
    g2439 <= gbuf187;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2440 <= 0;
  else
    g2440 <= g11582;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2441 <= 0;
  else
    g2441 <= gbuf188;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2442 <= 0;
  else
    g2442 <= g11583;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2443 <= 0;
  else
    g2443 <= gbuf189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2447 <= 0;
  else
    g2447 <= g11584;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2454 <= 0;
  else
    g2454 <= gbuf190;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2455 <= 0;
  else
    g2455 <= g11585;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2456 <= 0;
  else
    g2456 <= gbuf191;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2457 <= 0;
  else
    g2457 <= g11586;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2458 <= 0;
  else
    g2458 <= gbuf192;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2462 <= 0;
  else
    g2462 <= g11587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2469 <= 0;
  else
    g2469 <= gbuf193;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2470 <= 0;
  else
    g2470 <= g11588;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2471 <= 0;
  else
    g2471 <= gbuf194;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2472 <= 0;
  else
    g2472 <= g11589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2399 <= 0;
  else
    g2399 <= gbuf195;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2400 <= 0;
  else
    g2400 <= g13456;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2406 <= 0;
  else
    g2406 <= gbuf196;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2412 <= 0;
  else
    g2412 <= gbuf197;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2619 <= 0;
  else
    g2619 <= g13467;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2625 <= 0;
  else
    g2625 <= gbuf198;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2624 <= 0;
  else
    g2624 <= gbuf199;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2628 <= 0;
  else
    g2628 <= g23274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2631 <= 0;
  else
    g2631 <= g20568;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2584 <= 0;
  else
    g2584 <= g20569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2587 <= 0;
  else
    g2587 <= g16473;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2597 <= 0;
  else
    g2597 <= gbuf200;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2598 <= 0;
  else
    g2598 <= gbuf201;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2638 <= 0;
  else
    g2638 <= g11593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2643 <= 0;
  else
    g2643 <= gbuf202;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2644 <= 0;
  else
    g2644 <= g11596;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2645 <= 0;
  else
    g2645 <= gbuf203;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2646 <= 0;
  else
    g2646 <= g11597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2647 <= 0;
  else
    g2647 <= gbuf204;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2648 <= 0;
  else
    g2648 <= g11598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2639 <= 0;
  else
    g2639 <= gbuf205;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2640 <= 0;
  else
    g2640 <= g11594;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2641 <= 0;
  else
    g2641 <= gbuf206;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2642 <= 0;
  else
    g2642 <= g11595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2564 <= 0;
  else
    g2564 <= gbuf207;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2549 <= 0;
  else
    g2549 <= g13457;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2556 <= 0;
  else
    g2556 <= gbuf208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2560 <= 0;
  else
    g2560 <= gbuf209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2561 <= 0;
  else
    g2561 <= g24415;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2562 <= 0;
  else
    g2562 <= g24416;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2563 <= 0;
  else
    g2563 <= g24417;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2530 <= 0;
  else
    g2530 <= g25172;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2533 <= 0;
  else
    g2533 <= g25164;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2536 <= 0;
  else
    g2536 <= g25165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2552 <= 0;
  else
    g2552 <= g25169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2553 <= 0;
  else
    g2553 <= g25170;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2554 <= 0;
  else
    g2554 <= g25171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2555 <= 0;
  else
    g2555 <= g24412;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2559 <= 0;
  else
    g2559 <= g24413;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2539 <= 0;
  else
    g2539 <= g24414;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2540 <= 0;
  else
    g2540 <= g25166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2543 <= 0;
  else
    g2543 <= g25167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2546 <= 0;
  else
    g2546 <= g25168;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2602 <= 0;
  else
    g2602 <= g16474;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2609 <= 0;
  else
    g2609 <= gbuf210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2616 <= 0;
  else
    g2616 <= gbuf211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2617 <= 0;
  else
    g2617 <= g19057;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2618 <= 0;
  else
    g2618 <= gbuf212;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2622 <= 0;
  else
    g2622 <= g30325;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2623 <= 0;
  else
    g2623 <= g19058;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2574 <= 0;
  else
    g2574 <= gbuf213;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2632 <= 0;
  else
    g2632 <= g19059;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2633 <= 0;
  else
    g2633 <= gbuf214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2650 <= 0;
  else
    g2650 <= g28297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2651 <= 0;
  else
    g2651 <= g28298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2649 <= 0;
  else
    g2649 <= g28299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2653 <= 0;
  else
    g2653 <= g28300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2654 <= 0;
  else
    g2654 <= g28301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2652 <= 0;
  else
    g2652 <= g28302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2656 <= 0;
  else
    g2656 <= g28303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2657 <= 0;
  else
    g2657 <= g28304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2655 <= 0;
  else
    g2655 <= g28305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2659 <= 0;
  else
    g2659 <= g28306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2660 <= 0;
  else
    g2660 <= g28307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2658 <= 0;
  else
    g2658 <= g28308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2661 <= 0;
  else
    g2661 <= g26012;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2664 <= 0;
  else
    g2664 <= g26013;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2667 <= 0;
  else
    g2667 <= g26014;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2670 <= 0;
  else
    g2670 <= g26015;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2673 <= 0;
  else
    g2673 <= g26016;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2676 <= 0;
  else
    g2676 <= g26017;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2688 <= 0;
  else
    g2688 <= g29159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2691 <= 0;
  else
    g2691 <= g29160;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2694 <= 0;
  else
    g2694 <= g29161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2679 <= 0;
  else
    g2679 <= g29156;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2682 <= 0;
  else
    g2682 <= g29157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2685 <= 0;
  else
    g2685 <= g29158;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2565 <= 0;
  else
    g2565 <= g27233;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2568 <= 0;
  else
    g2568 <= g27234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2571 <= 0;
  else
    g2571 <= g27235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2580 <= 0;
  else
    g2580 <= g8311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2581 <= 0;
  else
    g2581 <= g24418;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2582 <= 0;
  else
    g2582 <= g19053;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2583 <= 0;
  else
    g2583 <= g19054;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2588 <= 0;
  else
    g2588 <= g19055;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2589 <= 0;
  else
    g2589 <= g19056;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2590 <= 0;
  else
    g2590 <= g30324;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2591 <= 0;
  else
    g2591 <= g30323;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2592 <= 0;
  else
    g2592 <= g30322;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2593 <= 0;
  else
    g2593 <= g30321;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2594 <= 0;
  else
    g2594 <= g30320;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2599 <= 0;
  else
    g2599 <= gbuf215;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2603 <= 0;
  else
    g2603 <= g13458;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2604 <= 0;
  else
    g2604 <= g13459;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2605 <= 0;
  else
    g2605 <= g13460;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2606 <= 0;
  else
    g2606 <= g13461;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2607 <= 0;
  else
    g2607 <= g13462;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2608 <= 0;
  else
    g2608 <= g13463;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2610 <= 0;
  else
    g2610 <= g13464;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2611 <= 0;
  else
    g2611 <= g13465;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2612 <= 0;
  else
    g2612 <= g26011;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2615 <= 0;
  else
    g2615 <= g13466;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2697 <= 0;
  else
    g2697 <= g13468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2700 <= 0;
  else
    g2700 <= gbuf216;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2703 <= 0;
  else
    g2703 <= gbuf217;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2704 <= 0;
  else
    g2704 <= g20570;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2733 <= 0;
  else
    g2733 <= g21946;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2714 <= 0;
  else
    g2714 <= g23275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2707 <= 0;
  else
    g2707 <= g24419;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2727 <= 0;
  else
    g2727 <= g25173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2720 <= 0;
  else
    g2720 <= g26018;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2734 <= 0;
  else
    g2734 <= g26742;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2746 <= 0;
  else
    g2746 <= g27236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2740 <= 0;
  else
    g2740 <= g27714;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2753 <= 0;
  else
    g2753 <= g28309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2760 <= 0;
  else
    g2760 <= g28692;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2766 <= 0;
  else
    g2766 <= g29162;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2773 <= 0;
  else
    g2773 <= g23276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2774 <= 0;
  else
    g2774 <= g23277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2772 <= 0;
  else
    g2772 <= g23278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2776 <= 0;
  else
    g2776 <= g23279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2777 <= 0;
  else
    g2777 <= g23280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2775 <= 0;
  else
    g2775 <= g23281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2779 <= 0;
  else
    g2779 <= g23282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2780 <= 0;
  else
    g2780 <= g23283;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2778 <= 0;
  else
    g2778 <= g23284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2782 <= 0;
  else
    g2782 <= g23285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2783 <= 0;
  else
    g2783 <= g23286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2781 <= 0;
  else
    g2781 <= g23287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2785 <= 0;
  else
    g2785 <= g23288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2786 <= 0;
  else
    g2786 <= g23289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2784 <= 0;
  else
    g2784 <= g23290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2788 <= 0;
  else
    g2788 <= g23291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2789 <= 0;
  else
    g2789 <= g23292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2787 <= 0;
  else
    g2787 <= g23293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2791 <= 0;
  else
    g2791 <= g23294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2792 <= 0;
  else
    g2792 <= g23295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2790 <= 0;
  else
    g2790 <= g23296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2794 <= 0;
  else
    g2794 <= g23297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2795 <= 0;
  else
    g2795 <= g23298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2793 <= 0;
  else
    g2793 <= g23299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2797 <= 0;
  else
    g2797 <= g23300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2798 <= 0;
  else
    g2798 <= g23301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2796 <= 0;
  else
    g2796 <= g23302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2800 <= 0;
  else
    g2800 <= g23303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2801 <= 0;
  else
    g2801 <= g23304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2799 <= 0;
  else
    g2799 <= g23305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2803 <= 0;
  else
    g2803 <= g23306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2804 <= 0;
  else
    g2804 <= g23307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2802 <= 0;
  else
    g2802 <= g23308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2806 <= 0;
  else
    g2806 <= g23309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2807 <= 0;
  else
    g2807 <= g23310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2805 <= 0;
  else
    g2805 <= g23311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2809 <= 0;
  else
    g2809 <= g26743;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2810 <= 0;
  else
    g2810 <= g26744;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2808 <= 0;
  else
    g2808 <= g26745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2812 <= 0;
  else
    g2812 <= g24420;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2813 <= 0;
  else
    g2813 <= g24421;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2811 <= 0;
  else
    g2811 <= g24422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3054 <= 0;
  else
    g3054 <= g23317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3079 <= 0;
  else
    g3079 <= g23318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3080 <= 0;
  else
    g3080 <= g21965;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3043 <= 0;
  else
    g3043 <= g29453;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3044 <= 0;
  else
    g3044 <= g29454;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3045 <= 0;
  else
    g3045 <= g29455;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3046 <= 0;
  else
    g3046 <= g29456;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3047 <= 0;
  else
    g3047 <= g29457;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3048 <= 0;
  else
    g3048 <= g29458;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3049 <= 0;
  else
    g3049 <= g29459;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3050 <= 0;
  else
    g3050 <= g29460;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3051 <= 0;
  else
    g3051 <= g29655;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3052 <= 0;
  else
    g3052 <= g29972;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3053 <= 0;
  else
    g3053 <= g29973;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3055 <= 0;
  else
    g3055 <= g29974;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3056 <= 0;
  else
    g3056 <= g29975;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3057 <= 0;
  else
    g3057 <= g29976;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3058 <= 0;
  else
    g3058 <= g29977;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3059 <= 0;
  else
    g3059 <= g29978;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3060 <= 0;
  else
    g3060 <= g29979;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3061 <= 0;
  else
    g3061 <= g30119;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3062 <= 0;
  else
    g3062 <= g30908;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3063 <= 0;
  else
    g3063 <= g30909;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3064 <= 0;
  else
    g3064 <= g30910;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3065 <= 0;
  else
    g3065 <= g30911;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3066 <= 0;
  else
    g3066 <= g30912;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3067 <= 0;
  else
    g3067 <= g30913;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3068 <= 0;
  else
    g3068 <= g30914;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3069 <= 0;
  else
    g3069 <= g30915;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3070 <= 0;
  else
    g3070 <= g30940;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3071 <= 0;
  else
    g3071 <= g30980;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3072 <= 0;
  else
    g3072 <= g30981;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3073 <= 0;
  else
    g3073 <= g30982;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3074 <= 0;
  else
    g3074 <= g30983;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3075 <= 0;
  else
    g3075 <= g30984;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3076 <= 0;
  else
    g3076 <= g30985;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3077 <= 0;
  else
    g3077 <= g30986;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3078 <= 0;
  else
    g3078 <= g30987;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2997 <= 0;
  else
    g2997 <= g30989;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2993 <= 0;
  else
    g2993 <= g26748;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2998 <= 0;
  else
    g2998 <= g27238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3006 <= 0;
  else
    g3006 <= g25177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3002 <= 0;
  else
    g3002 <= g26021;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3013 <= 0;
  else
    g3013 <= g26750;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3010 <= 0;
  else
    g3010 <= g27239;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3024 <= 0;
  else
    g3024 <= g27716;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3018 <= 0;
  else
    g3018 <= g24425;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3028 <= 0;
  else
    g3028 <= g25176;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3036 <= 0;
  else
    g3036 <= g26022;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3032 <= 0;
  else
    g3032 <= g26749;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3040 <= 0;
  else
    g3040 <= g16497;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2986 <= 0;
  else
    g2986 <= gbuf218;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2987 <= 0;
  else
    g2987 <= g16495;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g48 <= 0;
  else
    g48 <= g20595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g45 <= 0;
  else
    g45 <= g20596;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g42 <= 0;
  else
    g42 <= g20597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g39 <= 0;
  else
    g39 <= g20598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g27 <= 0;
  else
    g27 <= g20599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g30 <= 0;
  else
    g30 <= g20600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g33 <= 0;
  else
    g33 <= g20601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g36 <= 0;
  else
    g36 <= g20602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3083 <= 0;
  else
    g3083 <= g20603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g26 <= 0;
  else
    g26 <= g20604;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2992 <= 0;
  else
    g2992 <= g21966;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g23 <= 0;
  else
    g23 <= g20605;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g20 <= 0;
  else
    g20 <= g20606;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g17 <= 0;
  else
    g17 <= g20607;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g11 <= 0;
  else
    g11 <= g20608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g14 <= 0;
  else
    g14 <= g20589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5 <= 0;
  else
    g5 <= g20590;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g8 <= 0;
  else
    g8 <= g20591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2 <= 0;
  else
    g2 <= g20592;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2990 <= 0;
  else
    g2990 <= g20593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2991 <= 0;
  else
    g2991 <= g21964;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1 <= 0;
  else
    g1 <= g20594;
assign g18281 = ((~g14263));
assign g20592 = ((~II27101));
assign g29827 = (g29741&g22356);
assign g16081 = (g3304&g11783);
assign g24124 = ((~g22464));
assign g17318 = ((~II23406));
assign g29394 = ((~g29050));
assign II30149 = ((~g22736));
assign g13447 = ((~II20640));
assign g30503 = ((~g14213)&(~g30223));
assign g22225 = ((~II28789));
assign II39056 = ((~g29554));
assign g24850 = ((~g23464));
assign g23625 = (g22880&g20388);
assign II22919 = ((~g13945))|((~II22917));
assign g10306 = (g7162&g4665);
assign g17674 = (g4520&g15343);
assign g13491 = (g6028&g12221);
assign g28911 = ((~II37880));
assign g14745 = ((~II21289));
assign g28845 = ((~II37823))|((~II37824));
assign g30086 = (g29835&g11108);
assign g24831 = (g24100&g20401);
assign g24362 = ((~II31760));
assign g8508 = (g3566&g1627);
assign g6136 = ((~g672));
assign II14712 = ((~g138));
assign g30484 = (g30191&g11367);
assign g10300 = (g6945&g1257);
assign II37128 = ((~g28106));
assign II14615 = ((~g1842));
assign g11145 = ((~II18061));
assign g29928 = ((~g29673)&(~g22367));
assign II30754 = ((~g22074));
assign g26774 = (g26472&g19299);
assign II20550 = ((~g13267));
assign g27059 = (g23349&g26625);
assign g26797 = (g26148&g16659);
assign g30797 = ((~II40647));
assign g16015 = (g12013&g10859);
assign g20649 = ((~II27240));
assign g26716 = ((~II34755));
assign g6426 = ((~g1922));
assign g10764 = (g3834&g5391);
assign g26734 = ((~II34809));
assign g8932 = (g3494&g1183);
assign II32535 = ((~g23407));
assign g22800 = ((~II29582));
assign II29448 = ((~g20996));
assign g13576 = ((~g11650));
assign g24396 = ((~II31862));
assign g19524 = ((~g16924));
assign g6045 = ((~g2282));
assign II25037 = ((~g14071));
assign II36234 = ((~g27667));
assign II18509 = ((~g8770));
assign g30716 = ((~II40438));
assign g24600 = ((~II32184));
assign g25379 = ((~g24893));
assign II32323 = ((~g17927))|((~g23982));
assign g5845 = (g2412&g2428);
assign II28792 = ((~g21880));
assign II16965 = ((~g4734))|((~g4452));
assign g22712 = ((~II29392));
assign g20454 = ((~g17788));
assign g3250 = ((~II13146));
assign g13626 = ((~g11697));
assign g22527 = ((~II29077));
assign II21908 = ((~g13082));
assign g28160 = ((~g27422));
assign g7600 = ((~g2908));
assign II35964 = ((~g26826));
assign II27335 = ((~g19420));
assign II21819 = ((~g11710));
assign g27547 = ((~II35937));
assign g24903 = ((~II32642));
assign II40137 = ((~g30494));
assign g21458 = ((~II28003));
assign g26632 = ((~g25749));
assign g17865 = ((~II23926));
assign g22719 = (g14222&g21577);
assign g21081 = ((~g19940)&(~g18329));
assign g8862 = ((~II16114));
assign g4136 = ((~g862));
assign g8938 = ((~II16234));
assign g5913 = ((~g2120));
assign g23609 = (g4082&g22503);
assign II29372 = ((~g20968));
assign g18644 = ((~II24764))|((~II24765));
assign g9034 = (g6751&g1251);
assign II29125 = ((~g21777));
assign g25907 = ((~g24940));
assign II18100 = ((~g7265));
assign g22735 = ((~II29445));
assign II32851 = ((~g23694));
assign g23150 = ((~II29903));
assign g15647 = ((~II21900));
assign g28840 = (g5913&g28500);
assign g22695 = ((~II29357));
assign g7521 = ((~g2200));
assign g29308 = ((~II38459));
assign II25855 = ((~g1453))|((~g18110));
assign g19900 = (g1365&g18946);
assign g10560 = ((~g8008));
assign g29740 = ((~g29583)&(~g1914));
assign g24742 = ((~g23971)&(~g22869));
assign g22314 = ((~g20783));
assign g21780 = ((~g20255))|((~g6838));
assign g12193 = ((~g10432)&(~g10493)&(~g10555));
assign II22282 = ((~g2962))|((~g13348));
assign g25200 = ((~g24965))|((~g3306));
assign g22036 = (g21104&g21095&g21084&II28582);
assign g29098 = ((~II38085));
assign II34017 = ((~g25887));
assign II25857 = ((~g18110))|((~II25855));
assign g19765 = (g660&g18870);
assign II32695 = ((~g23858))|((~g14280));
assign II18314 = ((~g6369));
assign g17694 = (g7227&g16061);
assign II21793 = ((~g13123));
assign II25820 = ((~g1448))|((~II25819));
assign II33686 = ((~g25070));
assign II17200 = ((~g7936));
assign g22220 = (g21690&g12091);
assign g29295 = ((~g28823));
assign II34818 = ((~g26281));
assign g23556 = ((~II30614));
assign II29522 = ((~g21022));
assign g28186 = ((~g27535));
assign II36311 = ((~g27426));
assign II20514 = ((~g11769));
assign gbuf3 = (g2864);
assign g9635 = (g6232&g3937);
assign II22527 = ((~g13469));
assign g28168 = ((~g27459));
assign g10783 = ((~g7228));
assign g23276 = ((~II30281));
assign g28773 = ((~g15234)&(~g28465));
assign g28619 = ((~g28075));
assign g8106 = ((~II15369));
assign g29301 = ((~g28829));
assign g10230 = ((~II17200));
assign g19449 = (g16884&g14797&g14776);
assign g21375 = (g9342&g20374);
assign g17729 = ((~II23807))|((~II23808));
assign II40101 = ((~g30326));
assign g23536 = (g5963&g22829);
assign g27065 = ((~g24945)&(~g26029));
assign g14327 = (g7760&g12996);
assign II40832 = ((~g30811));
assign g21615 = ((~g16567)&(~g19957));
assign g10495 = (g6486&g614);
assign g27481 = ((~g27182)&(~g25980));
assign g19638 = (g4058&g17413);
assign g10186 = (g3013&g7466&g3024&II17156);
assign II17730 = ((~g7083));
assign g30816 = ((~II40700));
assign g29873 = ((~g29680));
assign g22625 = ((~g21113));
assign g6015 = ((~II14478));
assign g20573 = ((~II27044));
assign II26642 = ((~g17746));
assign g15809 = ((~g12657))|((~g6574));
assign g23984 = ((~II31226));
assign g4939 = ((~g1417));
assign II29656 = ((~g21070));
assign II18136 = ((~g5668));
assign g21135 = ((~g20114)&(~g20137)&(~g20160));
assign II40209 = ((~g30459));
assign g18334 = ((~II24346));
assign g8885 = ((~II16153));
assign g16039 = ((~g12756));
assign g21117 = ((~g20089)&(~g20110)&(~g20133));
assign g19028 = ((~II25147));
assign g14764 = ((~g11791));
assign g11650 = ((~g9080)&(~g9096)&(~g9105));
assign g22269 = ((~g21735)&(~g20044));
assign g6101 = ((~II14618));
assign g23183 = ((~II30002));
assign g24906 = (g18886&g23879);
assign g20420 = ((~g17637));
assign g29336 = (g29045&g29023);
assign g30376 = ((~II39933));
assign g28925 = ((~II37894));
assign g30833 = ((~II40751));
assign g8123 = ((~g144));
assign g4854 = ((~g2210));
assign g9109 = (g3774&g7724);
assign g25630 = ((~g24478));
assign g11565 = ((~II18671));
assign g16045 = (g12013&g10892);
assign g12868 = ((~II19929));
assign II15882 = ((~g3878));
assign II29145 = ((~g20891));
assign g4919 = ((~g1261));
assign II38178 = ((~g29098));
assign g25413 = ((~g24945));
assign II14489 = ((~g1496));
assign g30608 = ((~g30412)&(~g2605));
assign g16066 = (g12071&g10912);
assign g8817 = ((~II16031));
assign II23667 = ((~g15866));
assign g11907 = ((~g9927)&(~g10063)&(~g10154));
assign II21674 = ((~g11698));
assign g18465 = ((~II24501))|((~II24502));
assign II29399 = ((~g20977));
assign g23297 = ((~II30344));
assign g17652 = (g4480&g15326);
assign g11584 = ((~II18728));
assign g18048 = ((~g14053));
assign II23645 = ((~g13537));
assign g23313 = ((~II30392));
assign g13413 = ((~II20538));
assign g8704 = (g6643&g7996);
assign g13171 = ((~g8723)&(~g8755)&(~g8774));
assign g14158 = ((~g11974));
assign g22284 = ((~g21757)&(~g20081));
assign g15520 = (g8172&g12844);
assign II36379 = ((~g27682));
assign II33596 = ((~g24446));
assign g21876 = ((~g19792));
assign g10270 = (g7488&g4581);
assign II17919 = ((~g7976));
assign II19794 = ((~g10676));
assign g6142 = ((~g679));
assign II36993 = ((~g28034));
assign g30219 = (g30036&g8980);
assign II36690 = ((~g27319));
assign g28052 = ((~II36609));
assign g5989 = ((~g1576));
assign g19903 = (g2046&g18948);
assign g29575 = (g28813&g29402);
assign II40706 = ((~g30650));
assign g7264 = ((~II14942));
assign g5363 = ((~g3107));
assign g12921 = ((~g8958));
assign g13642 = (g6221&g12498);
assign g20790 = ((~II27379));
assign g3931 = ((~g171));
assign g5185 = ((~g1982));
assign g15179 = ((~II21476));
assign g27523 = ((~II35893));
assign II20526 = ((~g12519));
assign g11900 = ((~g11151));
assign II36601 = ((~g27295));
assign g29151 = ((~II38196));
assign g17136 = ((~g14768));
assign g10217 = (g3522&g4517);
assign g23051 = ((~g21121)&(~g21153));
assign II21313 = ((~g11743));
assign g25232 = ((~g24781)&(~g23600));
assign g10117 = (g6369&g4363);
assign II29675 = ((~g21075));
assign II20476 = ((~g9027));
assign g20273 = ((~g18795));
assign II23207 = ((~g9595))|((~g13867));
assign g30946 = (g30930&g20757);
assign g19156 = ((~II25351));
assign II34722 = ((~g26216));
assign g22142 = ((~g21402)&(~g19728));
assign g29246 = ((~II38345));
assign g15593 = (g7897&g13244);
assign g28361 = ((~g15729)&(~g28104));
assign g16392 = (g5940&g12052);
assign g5935 = ((~g948));
assign g27479 = ((~II35821));
assign g28059 = ((~g26034)&(~g27248));
assign g15148 = ((~II21461));
assign II38339 = ((~g29120));
assign II35028 = ((~g26513));
assign g30646 = ((~g16241)&(~g30445));
assign II35473 = ((~g27156));
assign g30764 = (g30628&g20837);
assign g22313 = ((~g20780));
assign g11811 = ((~g9606)&(~g9725)&(~g9809));
assign g20462 = ((~g17850));
assign g18994 = (g14895&g13657&g13677&g13706);
assign g14143 = (g8026&g12965);
assign g15989 = ((~II22163));
assign g20953 = ((~g19752)&(~g17695));
assign II29694 = ((~g21081));
assign g30469 = (g30159&g11281);
assign g24796 = (g12876&g24147);
assign g21020 = ((~g19852)&(~g17948));
assign g30333 = (g30191&g8341);
assign II31769 = ((~g23746));
assign g12599 = ((~g8763));
assign g26277 = ((~II34233));
assign g21550 = ((~II28080));
assign g30882 = ((~II40898));
assign g24519 = ((~g15459)&(~g23855));
assign g18389 = ((~II24408))|((~II24409));
assign g15210 = ((~g11840));
assign g30302 = ((~g13513)&(~g30003));
assign g27138 = ((~g26223));
assign g10400 = (g7230&g4845);
assign II37665 = ((~g28458));
assign II37488 = ((~g27765));
assign II21249 = ((~g11600));
assign g26301 = (g25258&g17749);
assign II40288 = ((~g30455));
assign g27184 = ((~g26085)&(~g25371));
assign g22638 = (g14001&g21498);
assign g8678 = ((~II15876));
assign II19542 = ((~g10574));
assign g20753 = ((~g20255))|((~g3722));
assign g4699 = ((~g2091));
assign g12804 = ((~II19865));
assign g20496 = ((~g18258));
assign g10405 = (g5556&g4865);
assign g29957 = (g29772&g29005);
assign g22467 = ((~II29013));
assign g4168 = ((~g1558));
assign g28151 = ((~g27381));
assign g26806 = ((~g15197)&(~g26244));
assign g4930 = ((~g1399));
assign II22924 = ((~g15118))|((~g14091));
assign g4720 = ((~g2498));
assign g19314 = ((~II25672))|((~II25673));
assign g12179 = ((~g10405)&(~g10468)&(~g10527));
assign II24539 = ((~g15118))|((~II24537));
assign g24446 = ((~g23433)&(~g22907));
assign g12485 = ((~II19667));
assign g24565 = (g20007&g18240&g23424);
assign II22845 = ((~g13579));
assign g29362 = ((~g28883));
assign g16881 = ((~II22860));
assign II39324 = ((~g29721))|((~II39323));
assign g28344 = ((~g15526)&(~g28027));
assign g30746 = ((~II40518));
assign II28494 = ((~g21358));
assign II31772 = ((~g23793));
assign g13194 = ((~g8784)&(~g8801)&(~g8816));
assign g21524 = ((~II28057));
assign g9582 = (g6369&g8215);
assign g10099 = ((~g7700));
assign g26480 = ((~II34444));
assign g24149 = ((~g22523));
assign g22246 = ((~g20659));
assign g25279 = ((~g24921)&(~g18140));
assign g30491 = ((~II40071));
assign g13656 = (g12776&g8640);
assign g15720 = ((~g12565))|((~g6232));
assign g7962 = ((~g1161));
assign g19843 = (g17741&g18190&II26285);
assign g26606 = ((~g25664));
assign g24069 = ((~g22922))|((~g14609));
assign g5305 = ((~g1997));
assign II13962 = ((~g2421));
assign II33858 = ((~g25179));
assign II32453 = ((~g24056))|((~II32451));
assign g17637 = ((~II23725));
assign g17252 = ((~II23338));
assign g26448 = ((~II34411));
assign g17704 = ((~II23788));
assign g17090 = (g7349&g15602);
assign g14114 = (g7718&g12951);
assign g13047 = ((~g9676))|((~g6980));
assign II18232 = ((~g6519));
assign g15867 = ((~g12611))|((~g6369));
assign g24427 = (g17086&g24134&g13626);
assign II17373 = ((~g3900));
assign g16345 = (g5897&g11971);
assign g16179 = ((~g12901));
assign II23894 = ((~g14177))|((~II23893));
assign II40218 = ((~g30335));
assign g5971 = ((~g2142));
assign g11731 = ((~g9968))|((~g3834));
assign g12041 = ((~g11370));
assign g11169 = ((~II18085));
assign g4702 = ((~g2109));
assign g13138 = ((~g9968))|((~g7426));
assign g25781 = ((~g24736)&(~g24523));
assign g10201 = (g3366&g4480);
assign g8556 = (g6838&g2270);
assign g29948 = (g29775&g28916);
assign g12122 = ((~g11478));
assign g4064 = ((~g1550));
assign g20836 = (g5829&g19125);
assign g26045 = ((~g25553)&(~g24885));
assign g8250 = ((~g2833));
assign g19312 = (g16924)|(g16578)|(g16529);
assign g20789 = ((~g19177)&(~g10340));
assign g16991 = (g7484&g15307);
assign g20614 = ((~II27167));
assign g10453 = (g5512&g4951);
assign II22900 = ((~g15022))|((~g14000));
assign II35000 = ((~g26336));
assign g22117 = ((~g21375)&(~g19679));
assign g30228 = ((~II39690))|((~II39691));
assign II33278 = ((~g25088));
assign g18803 = ((~g13704)&(~g11885));
assign II17992 = ((~g6314));
assign g18531 = ((~II24587))|((~II24588));
assign g7856 = ((~g3045));
assign g8257 = ((~g3201));
assign g11344 = ((~II18298));
assign g30245 = ((~g16074)&(~g30077));
assign II39541 = ((~g29913))|((~II39539));
assign g24300 = ((~II31574));
assign g23917 = (g7545&g23088);
assign g17954 = ((~g13992));
assign g27575 = ((~g26774)&(~g19107));
assign II33828 = ((~g25336));
assign g26357 = (g4882&g25634);
assign II34980 = ((~g26458));
assign g16767 = ((~II22759));
assign g16788 = ((~II22771));
assign g16446 = ((~g12611))|((~g3410));
assign g11506 = ((~II18494));
assign g27693 = ((~II36090));
assign II26726 = (g18735&g18765&g16266);
assign g26667 = ((~g25351)&(~g17149));
assign II16270 = ((~g5418));
assign g30689 = ((~g13486)&(~g30351));
assign g10328 = (g3774&g2498);
assign g5815 = ((~g991));
assign g25106 = ((~g24009))|((~g2059));
assign II28169 = ((~g19987));
assign g29485 = (g21508&g29290);
assign g9289 = ((~g5379));
assign II26440 = (g18603&g18555&g18504);
assign g13477 = (g6016&g12191);
assign g27401 = ((~II35741));
assign II27228 = ((~g19390));
assign g17901 = (g4902&g15531);
assign g12217 = ((~g10465)&(~g10526)&(~g10588));
assign g22276 = ((~g20714));
assign II20592 = ((~g11651));
assign g13366 = ((~II20455));
assign II21563 = ((~g13051));
assign g19668 = (g1339&g18827);
assign II30823 = ((~g21972));
assign g27756 = ((~g25410))|((~g27471));
assign g11045 = ((~II17960));
assign g7646 = ((~g318));
assign g5210 = ((~g2654));
assign g30986 = ((~II41132));
assign g24003 = ((~g22852))|((~g14537));
assign g26416 = (g5084&g25741);
assign g17143 = (g7685&g14099);
assign g18954 = ((~g15704));
assign II27119 = ((~g19563));
assign g19023 = ((~II25132));
assign g15602 = ((~g12363));
assign II16203 = ((~g3878));
assign II38459 = ((~g28749));
assign g25032 = ((~g23694))|((~g6713));
assign g25946 = ((~g24553)&(~g24561));
assign g24088 = ((~II31310));
assign g30265 = ((~g16349)&(~g30099));
assign II29357 = ((~g20965));
assign g25131 = ((~II32871));
assign g5142 = ((~g447));
assign g11759 = ((~g9302)&(~g9365)&(~g9438));
assign g8159 = ((~g1866));
assign g7896 = ((~II15212))|((~II15213));
assign g29996 = (g29901&g8443);
assign g18286 = ((~g14268));
assign II24716 = ((~g14497))|((~g9941));
assign g20342 = ((~g17378));
assign II18617 = ((~g11169));
assign II18461 = ((~g10931));
assign g10373 = (g6713&g4772);
assign II35425 = ((~g26832));
assign g8293 = ((~II15505));
assign g15304 = (g4573&g13192);
assign II36420 = ((~g27253));
assign g18917 = ((~g15557));
assign g11745 = ((~g10892));
assign g18003 = ((~g14024));
assign g14371 = ((~g12098));
assign g30550 = ((~II40230));
assign II13158 = ((~g165));
assign g10969 = ((~II17866));
assign g23215 = ((~II30098));
assign g23563 = (g8218&g22431);
assign II19174 = ((~g9263));
assign II13775 = ((~g109));
assign II40200 = ((~g30377));
assign II19739 = ((~g10694));
assign II13984 = ((~g1772));
assign g29973 = ((~II39457));
assign g16108 = (g5667&g11802);
assign g30682 = ((~g16450)&(~g30333));
assign g30568 = ((~g30402));
assign II31496 = ((~g23570));
assign g8915 = ((~II16203));
assign g3398 = ((~II13176));
assign g24359 = ((~II31751));
assign g29257 = (g28863&g8901);
assign II22063 = ((~g12999))|((~II22062));
assign g12233 = ((~g10477)&(~g10537)&(~g10596));
assign II38617 = ((~g28903));
assign g27904 = (g13873&g27387);
assign II29442 = ((~g20994));
assign II40484 = ((~g30677));
assign g10332 = ((~II17294));
assign II31670 = ((~g23463));
assign g30344 = ((~II39859));
assign g19142 = (g17159&g16719);
assign g27133 = ((~g26105));
assign g26145 = ((~g6068)&(~g24183)&(~g25347));
assign II28594 = (g21167&g21147&g21134);
assign g30010 = ((~g29520)&(~g29942));
assign II16321 = ((~g5425));
assign g10007 = (g6314&g4205);
assign II32919 = ((~g24560));
assign II33633 = ((~g24524));
assign g30526 = ((~II40158));
assign g11550 = ((~II18626));
assign g24493 = ((~g23693)&(~g22614));
assign g26614 = ((~g25688));
assign II26960 = ((~g16884));
assign g9111 = (g5556&g7730);
assign g7676 = ((~g402));
assign II15256 = ((~g2950));
assign g30296 = ((~g13488)&(~g29993));
assign g27508 = ((~II35868));
assign g18884 = ((~g13469));
assign g13559 = ((~g12657))|((~g3566));
assign g24034 = ((~g22812))|((~g14252));
assign g10854 = ((~II17705));
assign II22783 = ((~g13572));
assign g10333 = ((~II17297));
assign g26469 = (g5249&g25827);
assign g5894 = ((~g186));
assign II25838 = ((~g88))|((~g17802));
assign g30403 = ((~g30004)&(~g30131));
assign g26206 = ((~II34124));
assign II18211 = ((~g6232));
assign g13098 = ((~g9534))|((~g6678));
assign g20133 = (g18170&g9505);
assign g10616 = (g7015&g5246);
assign g30288 = ((~g16454)&(~g29984));
assign g27422 = ((~II35762));
assign g6029 = ((~II14496));
assign II40605 = ((~g30610))|((~II40603));
assign II24292 = ((~g9203))|((~II24290));
assign g12340 = ((~II19507));
assign g25977 = (g24845&g12089);
assign g28337 = (g28002&g19448);
assign g29175 = (g29009&g20687);
assign g27317 = ((~g27059)&(~g26408));
assign g25627 = (g24505&g20477);
assign g29943 = ((~II39423));
assign II31784 = ((~g23863));
assign II25111 = ((~g18981));
assign g18656 = ((~g14776));
assign g24257 = (g14381)|(g22365);
assign g12505 = ((~g8646));
assign g19201 = (g18183)|(g18424);
assign II32159 = ((~g24226));
assign g5766 = ((~g990));
assign g28211 = ((~II36882));
assign g22657 = ((~II29277));
assign II39157 = ((~g29618));
assign g4283 = ((~g1808));
assign g20526 = ((~g18446));
assign g10165 = (g7358&g4412);
assign g23489 = ((~g22850))|((~g14529))|((~g10714));
assign g30779 = ((~II40604))|((~II40605));
assign II25606 = ((~g744))|((~II25605));
assign II34686 = ((~g26398));
assign II19412 = ((~g10486));
assign II18455 = ((~g11031));
assign g26872 = ((~II35053));
assign g16708 = ((~g14849));
assign II38807 = ((~g29356));
assign II23556 = ((~g15837));
assign g26826 = ((~g15508)&(~g26391));
assign g14309 = ((~g12057));
assign g19861 = (g2734&g18924);
assign g11108 = ((~II18022));
assign g13373 = ((~g10482));
assign g8640 = ((~II15830));
assign g20307 = (g13764&g16360&II26726);
assign g9919 = (g7162&g4147);
assign g14554 = ((~g12216));
assign g25261 = ((~g24861)&(~g23796));
assign g18811 = ((~g15136));
assign g25994 = ((~II33834));
assign g27298 = ((~g27032)&(~g26366));
assign g30159 = ((~g30016));
assign g8844 = ((~II16082));
assign g27946 = ((~II36411));
assign g17157 = ((~g13552));
assign g13022 = ((~g8566)&(~g8573)&(~g8576));
assign g29288 = ((~II38421));
assign g18653 = (g14811&g14910&g13687&g16254);
assign g27794 = ((~II36243));
assign II19759 = ((~g10714));
assign gbuf130 = (g1663);
assign II35413 = ((~g26876));
assign g16733 = ((~II22745));
assign II24131 = ((~g14107))|((~g9471));
assign g14060 = ((~g8605))|((~g12515));
assign II31889 = ((~g23845));
assign g19192 = (g18183)|(g18270);
assign g11022 = ((~II17933));
assign II16062 = ((~g3900));
assign g29641 = ((~II39041));
assign g26697 = ((~II34698));
assign g23595 = ((~II30689));
assign g17248 = ((~g16052)&(~g16072));
assign g6977 = ((~g1145));
assign g16074 = (g5646&g11782);
assign II18192 = ((~g7895))|((~II18190));
assign g29340 = ((~g28337)&(~g28722));
assign g25165 = ((~II32973));
assign g27590 = ((~g27144));
assign g21939 = ((~g20040));
assign g16484 = ((~II22554));
assign g26902 = ((~g25631))|((~g26283))|((~g25569));
assign g17219 = ((~g4671)&(~g14584));
assign g29478 = (g21580&g29277);
assign g13219 = ((~g9770));
assign g13226 = ((~g9876));
assign g19282 = (g16954&g14507&g14423);
assign g13420 = ((~II20559));
assign g25596 = ((~II33421));
assign g24237 = ((~g17081)&(~g22311));
assign g15251 = ((~II21534));
assign g22412 = ((~II28956));
assign g11324 = ((~II18274));
assign II15213 = ((~g2953))|((~II15211));
assign gbuf35 = (g288);
assign g21097 = (g19505&g14273&g16507);
assign g10729 = (g7426&g5375);
assign g27923 = (g4144&g27419);
assign II28019 = ((~g20025));
assign II15012 = ((~g2700));
assign g28220 = ((~II36909));
assign II19986 = ((~g8577));
assign II17889 = ((~g6314));
assign II32143 = ((~g24218));
assign II14195 = ((~g3212));
assign g19782 = (g4538&g17685);
assign g24846 = (g24109&g20426);
assign g21913 = (g4456&g20519);
assign II32189 = ((~g24243));
assign g27310 = ((~g27050)&(~g26392));
assign g28612 = ((~g28046));
assign II18545 = ((~g8630));
assign II26377 = (g18521&g14119&g14217);
assign II27927 = ((~g19957));
assign g23863 = ((~II31115));
assign II13578 = ((~g1481));
assign g23476 = (g18643&g22661);
assign II40091 = ((~g30266));
assign g18188 = ((~g14252));
assign g23289 = ((~II30320));
assign g15562 = (g5088&g13240);
assign g13251 = ((~g8868)&(~g8899)&(~g8932));
assign g28761 = ((~g28445)&(~g27936));
assign II37020 = ((~g27910));
assign II31056 = ((~g22164));
assign g19721 = (g2707&g18848);
assign gbuf211 = (g2609);
assign g10043 = (g6519&g4240);
assign g28524 = ((~II37467));
assign g10653 = ((~g8159));
assign g28903 = ((~g28660)&(~g13295));
assign g23941 = (g18526&g23098);
assign II31802 = ((~g23460));
assign II17140 = ((~g3806));
assign g7709 = ((~g1006));
assign g7950 = ((~g142));
assign II35856 = ((~g26809));
assign g21211 = ((~g19240)&(~g19230));
assign g28108 = ((~II36755));
assign g27252 = ((~g26963)&(~g26207));
assign g19720 = (g4301&g17551);
assign g8026 = ((~g3060));
assign g25833 = ((~II33673));
assign g23234 = ((~II30155));
assign II36486 = ((~g27507));
assign II27050 = ((~g19183));
assign g17597 = (g6977&g16039);
assign g20385 = ((~g17514));
assign II37599 = ((~g28553));
assign II36250 = ((~g27612));
assign g12005 = ((~g10174)&(~g10261)&(~g10328));
assign II40515 = ((~g30687));
assign g23974 = ((~g4632)&(~g13573)&(~g23025));
assign g17578 = (g4354&g15254);
assign g27772 = (g5680&g27465);
assign II37800 = ((~g28635));
assign g23433 = ((~g22726)&(~g21611));
assign g22980 = ((~g21794));
assign II37965 = ((~g28529));
assign g29181 = ((~g28850)&(~g28407));
assign g13428 = ((~II20583));
assign g17177 = ((~g14118))|((~g14041));
assign g24973 = ((~g23819));
assign g12157 = ((~g8347));
assign II33813 = ((~g25706));
assign g29093 = ((~II38074));
assign g22196 = (g21597&g21012);
assign II25445 = ((~g18968));
assign g16265 = (g5823&g11910);
assign g7610 = ((~g312));
assign g28177 = ((~g27510));
assign II32952 = ((~g24570));
assign g22750 = ((~II29484));
assign g19185 = ((~II25406));
assign II35548 = ((~g27116));
assign II34156 = ((~g25235));
assign g8490 = (g6369&g945);
assign II24005 = ((~g7548))|((~g15814));
assign g15118 = ((~g11807));
assign II37011 = ((~g28078));
assign g9426 = ((~g5543));
assign g20220 = (g18593&g9355);
assign II13239 = ((~g2704));
assign g19710 = (g1332&g18843);
assign g15747 = ((~II21995));
assign g29267 = ((~II38386));
assign g14059 = (g7697&g12934);
assign II36358 = ((~g27672));
assign II25089 = ((~g14991));
assign g25533 = ((~II33361));
assign II27014 = ((~g19151));
assign g24411 = ((~II31907));
assign II32892 = ((~g24582));
assign II41090 = ((~g30965));
assign g13498 = (g6033&g12251);
assign g26610 = ((~g25675));
assign II27008 = ((~g19175));
assign II24763 = ((~g6194))|((~g14573));
assign g17212 = ((~II23292));
assign g21609 = (g19084)|(g16954)|(g14423);
assign II41114 = ((~g30976));
assign g19226 = (g18147)|(g18231);
assign g22045 = ((~g21312)&(~g19572));
assign g23693 = (g17914&g23002);
assign g10463 = (g3678&g4973);
assign g13540 = ((~g12657))|((~g3566));
assign g15496 = ((~II21755));
assign II38151 = ((~g29082));
assign II18731 = ((~g8945));
assign g23077 = ((~g14577)&(~g14524)&(~g21182));
assign g15997 = ((~g12561));
assign II18001 = ((~g6643));
assign g9366 = (g6232&g8059);
assign g26572 = ((~g25557));
assign g13610 = ((~II20832));
assign g12689 = ((~g8798));
assign II32074 = ((~g23413));
assign II19466 = ((~g10631));
assign g23410 = ((~g23071));
assign g8434 = ((~II15636));
assign II23966 = ((~g14092))|((~g9248));
assign g18719 = ((~g13643)&(~g13656));
assign g12775 = ((~g8832));
assign g12424 = ((~g10962));
assign g9048 = (g3338&g489);
assign II38801 = ((~g29358));
assign II33482 = ((~g24454));
assign g18939 = ((~g15644));
assign g16351 = ((~g13036));
assign II19449 = ((~g10424));
assign II34830 = ((~g26349));
assign g23252 = ((~II30209));
assign g19289 = (g17029&g8580);
assign II23854 = ((~g15970));
assign II15629 = ((~g5837));
assign II34233 = ((~g25250));
assign g5829 = ((~g1686));
assign II35399 = ((~g26199));
assign g28804 = ((~II37765));
assign II16095 = ((~g6082));
assign g16426 = (g5969&g12103);
assign g19118 = ((~II25315));
assign II17837 = ((~g8031));
assign g21476 = (g9569&g20442);
assign g25067 = ((~g24249)&(~g17100));
assign II31484 = ((~g23568));
assign gbuf121 = (g1517);
assign g15843 = ((~g12565))|((~g6314));
assign g21306 = (g9187&g20298);
assign II33504 = ((~g25037));
assign g18726 = ((~g13645)&(~g11805));
assign g27692 = ((~II36087));
assign II39008 = ((~g29509));
assign II16918 = ((~g6751));
assign g25057 = ((~g23748))|((~g5512));
assign g8455 = ((~II15657));
assign g21032 = ((~g19870)&(~g17990));
assign g15889 = ((~g12611))|((~g6369));
assign g24014 = ((~II31244));
assign g28693 = ((~II37626));
assign g22204 = ((~g19939)&(~g21681));
assign II17750 = ((~g7157));
assign g20516 = ((~g18432));
assign g21746 = ((~g14378))|((~g15263))|((~g19902))|((~g19875));
assign II36705 = ((~g27323));
assign II38737 = ((~g29339));
assign g29005 = ((~II37968));
assign gbuf23 = (g135);
assign g30866 = ((~II40850));
assign g22869 = (g14596&g21700);
assign g11876 = ((~g11108));
assign g30521 = ((~II40143));
assign g28255 = ((~II37014));
assign g22576 = ((~g17111)&(~g21925));
assign g14703 = ((~II21271));
assign g19232 = (g18302)|(g18514);
assign g30677 = ((~g16421)&(~g30499));
assign II21708 = ((~g13081));
assign II34737 = ((~g26439));
assign g22147 = ((~g21413)&(~g19738));
assign g12847 = ((~g8882));
assign II21742 = ((~g13114));
assign g7869 = ((~g2959));
assign g20043 = ((~g18240));
assign g10102 = (g6314&g4332);
assign g11943 = ((~g11222));
assign g22179 = ((~g21481)&(~g19813));
assign g29833 = (g29725&g20813);
assign II38951 = ((~g29221));
assign gbuf76 = (g1092);
assign g10175 = (g5556&g4438);
assign g19828 = (g2734&g18905);
assign g7358 = ((~II14976));
assign g7193 = ((~g1491));
assign g20311 = ((~g17304));
assign g30026 = ((~g29560)&(~g29959));
assign g25667 = ((~II33491));
assign g30123 = (g30070&g20641);
assign g15603 = ((~g12366));
assign II25432 = ((~g18837));
assign g30593 = ((~g30412)&(~g2603));
assign g20693 = ((~g20228))|((~g3566));
assign g8531 = (g3254&g201);
assign g26154 = ((~g6068)&(~g24183)&(~g25329));
assign g19982 = (g17992&g17913&II26432);
assign II36321 = ((~g27627));
assign g11222 = ((~II18148));
assign g19490 = ((~g16761));
assign II22581 = ((~g14766));
assign g15388 = (g7834&g12769);
assign II40600 = ((~g30707));
assign g15810 = ((~g12657))|((~g6783));
assign g21751 = ((~II28272))|((~II28273));
assign g19245 = (g18395)|(g18578);
assign g22606 = (g2720&g21876);
assign II25500 = (g17058)|(g17030)|(g17016);
assign g4094 = ((~g3207));
assign g26118 = ((~II34012));
assign g11884 = ((~g11123));
assign II36063 = ((~g27463));
assign g27086 = (g23353&g26643);
assign g11767 = ((~g9366)&(~g9439)&(~g9518));
assign II19404 = ((~g10664));
assign g27702 = ((~II36117));
assign g25967 = ((~g24596)&(~g23512));
assign II29812 = ((~g21467));
assign g20895 = ((~g19633)&(~g17461));
assign g13400 = ((~g10545));
assign g22186 = ((~g21497)&(~g19837));
assign II34698 = ((~g26181));
assign g26441 = (g5170&g25784);
assign g30382 = ((~II39951));
assign g29638 = ((~II39032));
assign g27570 = (g24038&g27173);
assign g10880 = ((~II17743));
assign g15640 = (g5217&g13263);
assign II30026 = ((~g22586));
assign II18929 = ((~g10711));
assign g4611 = ((~g710));
assign g11989 = ((~g11297));
assign g10918 = ((~II17801));
assign g29911 = ((~II39324))|((~II39325));
assign g13432 = ((~II20595));
assign g22660 = (g14053&g21524);
assign g21226 = (g20242&g12426);
assign g20335 = ((~g17366));
assign g29515 = ((~II38875));
assign g10204 = (g6912&g4489);
assign g21268 = (g19641&g15065);
assign g11834 = ((~g11036));
assign g21970 = ((~g17182)&(~g21226));
assign g17416 = ((~II23504));
assign II31115 = ((~g22180));
assign g8620 = ((~II15806));
assign g22948 = ((~II29727));
assign g18735 = ((~g14922));
assign g21812 = (g16705&g19608&g14811);
assign g12265 = ((~g8452));
assign II20909 = ((~g13055));
assign g4307 = ((~g2252));
assign g21823 = (g20218)|(g20186)|(g18638)|(g19116);
assign g11237 = ((~II18163));
assign II33611 = ((~g25055));
assign g23064 = ((~g21612));
assign g30061 = ((~g29971)&(~g13493));
assign g24009 = ((~g23017)&(~g7259));
assign II37291 = ((~g28148));
assign g12978 = ((~g8529)&(~g8544)&(~g8557));
assign g7926 = ((~g3067));
assign g15723 = ((~g12611))|((~g6519));
assign g24824 = (g9857&g24165);
assign g27907 = ((~II36362));
assign g13853 = (g7580&g12689);
assign g26442 = ((~II34405));
assign g17630 = (g4314&g16042);
assign g23663 = ((~II30803));
assign g23459 = ((~II30493));
assign II26426 = ((~g16536));
assign g25758 = ((~II33589));
assign g24160 = ((~g22540));
assign g29661 = ((~g29576));
assign g15659 = ((~g11706));
assign g4395 = ((~g1543));
assign g11682 = ((~II18866));
assign II30350 = ((~g22901));
assign g19254 = (g16895&g14273&g14186);
assign g20053 = (g17720&g12875);
assign II40471 = ((~g30673));
assign g28242 = ((~II36975));
assign II40961 = ((~g30749));
assign g21846 = (g20249)|(g18648)|(II28369);
assign g21446 = (g9711&g20429);
assign g27119 = ((~g26367))|((~g6713));
assign II26195 = ((~g16853));
assign g14573 = ((~g12233));
assign g30670 = ((~g16389)&(~g30484));
assign g27435 = ((~g26777)&(~g25193));
assign g6309 = ((~g14));
assign g9758 = ((~g5618));
assign II14556 = ((~g1142));
assign g26753 = ((~II34866));
assign g10466 = (g3722&g4982);
assign g16479 = ((~II22539));
assign II23035 = ((~g9232))|((~II23034));
assign g13075 = ((~g9676))|((~g7162));
assign g18942 = ((~g13870)&(~g12273));
assign g16091 = ((~g12825));
assign g3984 = ((~g2222));
assign II14631 = ((~g2473));
assign g4115 = ((~g698));
assign g13356 = ((~II20441));
assign g25706 = ((~II33532));
assign II40164 = ((~g30446));
assign II14574 = ((~g1750));
assign g13816 = (g7530&g12596);
assign g23009 = ((~g21738)&(~g21107));
assign g22458 = ((~II29004));
assign g23854 = (g18265&g23049);
assign g10365 = (g3338&g593);
assign g20406 = ((~g17588));
assign g19971 = (g5327&g18355);
assign g28102 = ((~II36741));
assign g19803 = (g666&g18892);
assign II33182 = ((~g25056));
assign g22549 = ((~II29101));
assign II22316 = ((~g2934))|((~g13370));
assign g17556 = (g4201&g16027);
assign g5149 = ((~g617));
assign II37188 = ((~g27785));
assign g7538 = ((~g2536));
assign g28472 = (g18207&g27959);
assign g5888 = ((~g2615));
assign g13518 = ((~g12565))|((~g3254));
assign II40254 = ((~g30474));
assign g20292 = ((~g17265));
assign g17122 = (g7658&g14024);
assign g19808 = (g1358&g18897);
assign II39401 = ((~g29662));
assign g17042 = ((~g14691)&(~g14669)&(~g15890));
assign g25451 = ((~g16048)&(~g25102));
assign II17054 = ((~g7391));
assign g28466 = (g26131&g28170);
assign II19952 = ((~g8571));
assign II18444 = ((~g7391));
assign g23627 = ((~II30751));
assign II24587 = ((~g14596))|((~II24586));
assign g26835 = ((~II34974));
assign g15240 = ((~II21523));
assign II25580 = ((~g18281))|((~II25578));
assign II23478 = ((~g15844));
assign g22154 = ((~g21424)&(~g19756));
assign g15410 = (g4786&g13208);
assign g18850 = ((~g15314));
assign g26957 = ((~g26577));
assign II37885 = ((~g28556));
assign II23075 = ((~g9293))|((~II23074));
assign II37459 = ((~g27759));
assign II22917 = ((~g15096))|((~g13945));
assign II26574 = ((~g18325));
assign g19883 = (g4982&g17951);
assign g5326 = ((~g2873));
assign II18181 = ((~g5636));
assign II13232 = ((~g2624));
assign g30229 = ((~g30030));
assign g30963 = ((~g30957));
assign g24078 = ((~g22887))|((~g14408));
assign g29761 = ((~g28707)&(~g28711)&(~g29466));
assign g25405 = ((~g24933));
assign g28997 = (g28630&g9623);
assign II38119 = ((~g28420));
assign g26882 = ((~g25514)&(~g26301));
assign g11887 = ((~g11129));
assign II16303 = ((~g6713));
assign g9630 = (g3254&g3922);
assign g26240 = ((~g25968)&(~g13340));
assign II25311 = (g18744&g18772&g18815);
assign II37379 = ((~g28199));
assign g25110 = ((~g23867));
assign g6066 = ((~II14577));
assign g18183 = ((~II24179))|((~II24180));
assign g28381 = (g28157&g9815);
assign g21335 = (g9248&g20331);
assign g26821 = ((~g15424)&(~g26347));
assign g30756 = ((~II40542));
assign g9936 = ((~II16942));
assign II28000 = ((~g19167));
assign g30949 = (g30933&g20806);
assign g25022 = ((~g23694))|((~g6713));
assign g22705 = ((~II29375));
assign II32430 = ((~g17815))|((~g24052));
assign g29464 = (g29190&g8375);
assign II30374 = ((~g22775));
assign II16653 = ((~g5512));
assign II38821 = ((~g29313))|((~II38820));
assign g17878 = ((~g15830));
assign g10911 = ((~II17792));
assign II18677 = ((~g8908));
assign g16061 = ((~g12798));
assign II25655 = ((~g17937))|((~II25653));
assign g12645 = ((~g8785));
assign g21040 = ((~g19880)&(~g18036));
assign g5412 = ((~II13950));
assign g4409 = ((~g2078));
assign II30741 = ((~g22068));
assign g14882 = ((~II21337));
assign g29510 = ((~II38860));
assign g13280 = ((~II20339));
assign II22810 = ((~g14280));
assign g12328 = ((~g10641)&(~g10672)&(~g10690));
assign II20637 = ((~g11652));
assign II40098 = ((~g30491));
assign g16863 = ((~II22845));
assign g9766 = (g5438&g4017);
assign II28712 = ((~g21851));
assign g9160 = ((~g6170));
assign g24337 = ((~II31685));
assign g21298 = (g9356&g20286);
assign II36411 = ((~g27582));
assign g25019 = ((~g23923))|((~g6486));
assign g11672 = ((~g9534))|((~g3366));
assign g5400 = ((~II13916));
assign g17998 = ((~II24037))|((~II24038));
assign g27236 = ((~II35545));
assign g10586 = (g7358&g5190);
assign II27232 = ((~g19401));
assign g25239 = ((~g24796)&(~g23615));
assign g19597 = (g3922&g17342);
assign g20974 = ((~g19776)&(~g17754));
assign g17012 = ((~g14657)&(~g14642)&(~g15859));
assign g10599 = (g3834&g5227);
assign II22599 = ((~g14966));
assign g10475 = (g3834&g5009);
assign g12197 = ((~g8391));
assign g4237 = ((~g844));
assign g23052 = (g21800)|(g21788)|(g21844);
assign II29077 = ((~g20718));
assign g20157 = (g18415&g9287);
assign g15494 = (g4962&g13223);
assign II37334 = ((~g28194));
assign II38232 = ((~g29117));
assign g25655 = ((~II33479));
assign g15557 = ((~II21813));
assign g9257 = ((~II16511));
assign g23174 = ((~II29975));
assign g24180 = ((~g22629));
assign g26390 = (g25919&g9873);
assign II24205 = ((~g6568))|((~g14102));
assign II13173 = ((~g629));
assign g19932 = (g2917&g18166);
assign g23452 = ((~II30480));
assign II38725 = ((~g29327));
assign gbuf55 = (g564);
assign g24098 = ((~g22409));
assign II14149 = ((~g3231));
assign g13805 = ((~g12471));
assign g27697 = ((~II36102));
assign II25733 = ((~g18091))|((~II25731));
assign g22834 = ((~II29625));
assign g12172 = ((~g10400)&(~g10464)&(~g10525));
assign II19025 = ((~g9225));
assign g29431 = ((~II38674));
assign g12819 = ((~g9248)&(~g9203));
assign II38958 = ((~g29226));
assign II37578 = ((~g28432));
assign g22810 = ((~g16075)&(~g20842)&(~g21271));
assign II35821 = ((~g26804));
assign g15827 = ((~g12711))|((~g7085));
assign g13621 = ((~g12955))|((~g3678));
assign II14538 = ((~g369));
assign II23501 = ((~g15825));
assign g10935 = ((~II17828));
assign II35554 = ((~g27102));
assign g9442 = (g6232&g8135);
assign II38447 = ((~g28744));
assign II40784 = ((~g30813));
assign g26562 = ((~g25527));
assign II30598 = ((~g22027));
assign II19303 = ((~g9422));
assign g19042 = ((~II25189));
assign g17529 = (g4260&g15204);
assign g29226 = ((~g15374)&(~g28997));
assign g27315 = ((~g27057)&(~g26405));
assign g3238 = ((~II13110));
assign g24536 = ((~g23877)&(~g22745));
assign g22451 = ((~II28997));
assign II40227 = ((~g30350));
assign II20532 = ((~g13339));
assign g30937 = ((~II41035));
assign g27747 = ((~g27427)&(~g26973));
assign II38536 = ((~g28920));
assign g8341 = ((~II15543));
assign g27032 = (g22005&g26603);
assign g21354 = (g9264&g20352);
assign g10515 = (g3618&g5072);
assign g25253 = ((~g24826)&(~g23681));
assign g14230 = ((~II21127));
assign g23746 = ((~II30944));
assign g10649 = ((~g3398))|((~g6912));
assign g27466 = ((~g26915)&(~g24624));
assign g11669 = ((~g9099)&(~g9108)&(~g9115));
assign II16930 = (g5942&g4683&g4684&g5297);
assign g21330 = (g9150&g20329);
assign II28249 = ((~g19494))|((~II28247));
assign II23908 = ((~g14337));
assign g23579 = (g3963&g22461);
assign g22533 = ((~II29083));
assign g26686 = ((~II34665));
assign g26367 = (g25873)|(g25882);
assign II23191 = ((~g9507))|((~II23190));
assign g29192 = ((~g28954));
assign II29016 = ((~g21696));
assign g10255 = (g6838&g4558);
assign II36571 = ((~g27288));
assign g5907 = ((~g1618));
assign g5835 = ((~g2291));
assign II18402 = ((~g6713));
assign g24588 = ((~II32156));
assign II16726 = ((~g6085));
assign g29508 = ((~II38854));
assign g19206 = (g18053)|(g18319);
assign g7906 = ((~g488));
assign II15167 = ((~g2981))|((~g2874));
assign g26022 = ((~II33918));
assign g10396 = (g3678&g4833);
assign g28316 = ((~II37197));
assign II24474 = ((~g6184))|((~g14580));
assign II35410 = ((~g26872));
assign g12024 = ((~g11354));
assign II37137 = ((~g28117));
assign II21680 = ((~g13102));
assign g17021 = (g7592&g15438);
assign g27834 = ((~g27478)&(~g14630));
assign g30371 = ((~II39922));
assign g29220 = (g15296&g28779);
assign g23512 = (g5858&g22328);
assign g11515 = ((~II18521));
assign g22676 = ((~II29320));
assign g15516 = ((~II21775));
assign g28249 = ((~II36996));
assign II17294 = ((~g7936));
assign g20098 = (g18383)|(g18302)|(II26532);
assign II14647 = ((~g2543));
assign g15873 = ((~g11617)&(~g7562));
assign g16453 = (g5989&g12157);
assign g11051 = ((~II17966));
assign g24572 = ((~II32120));
assign II32422 = ((~g18155))|((~g24046));
assign g22685 = ((~II29339));
assign II16309 = ((~g5512));
assign II21952 = ((~g13132));
assign g26083 = ((~g25426)&(~g22319));
assign g10321 = (g7230&g4699);
assign g30854 = ((~II40814));
assign g11651 = ((~II18835));
assign g16986 = ((~II22925))|((~II22926));
assign g26768 = (g26440&g19280);
assign II34400 = ((~g25267));
assign g15688 = ((~II21939));
assign g17018 = (g7830&g15409);
assign g22915 = ((~g19491))|((~g20928));
assign II17895 = ((~g6448));
assign II30002 = ((~g22730));
assign g10679 = ((~g3554))|((~g7162));
assign II16190 = ((~g6118));
assign g19736 = (g4360&g17579);
assign g17755 = ((~II23830));
assign g13297 = ((~g10232));
assign g8354 = ((~II15556));
assign II40475 = ((~g30674));
assign g13482 = ((~g12657))|((~g3566));
assign g26428 = ((~II34385));
assign g24083 = ((~g22015)&(~g20836));
assign g26006 = ((~II33870));
assign g27279 = ((~g27007)&(~g26324));
assign II30908 = ((~g22123));
assign g29639 = ((~II39035));
assign g11188 = ((~II18107))|((~II18108));
assign g27251 = ((~g26958)&(~g26186));
assign II32492 = ((~g24067))|((~II32490));
assign g13469 = ((~II20706));
assign g20333 = ((~g13672)&(~g16859));
assign II23368 = ((~g16446));
assign g29436 = ((~II38689));
assign g17017 = (g7590&g15408);
assign g26062 = (g25947&g21113);
assign g28738 = ((~g14975)&(~g28433));
assign g21083 = ((~g19943)&(~g18333));
assign g22385 = ((~g21207))|((~g21266))|((~g21196));
assign II25672 = ((~g2160))|((~II25671));
assign II18575 = ((~g8845));
assign g25489 = (g24795)|(g16466);
assign g29781 = ((~g29481)&(~g29233));
assign g17282 = ((~II23368));
assign g25151 = ((~II32931));
assign g15990 = ((~g12886))|((~g6912));
assign II18082 = ((~g6574));
assign II41105 = ((~g30968));
assign II29291 = ((~g20940));
assign g29049 = ((~g9248))|((~g28540));
assign g8690 = ((~II15890));
assign g19018 = ((~II25117));
assign g28141 = ((~g27576));
assign g19542 = (g16974)|(g16797)|(g16743);
assign II31724 = ((~g23581));
assign g21859 = ((~g18030))|((~g19195))|((~g19204));
assign g6421 = ((~g1326));
assign g28421 = ((~g16068)&(~g28176));
assign g17682 = ((~II23766));
assign g10630 = (g5556&g5266);
assign g24037 = ((~g22887))|((~g14592));
assign g30968 = ((~g30960));
assign g25770 = ((~II33603));
assign II32660 = ((~g18038))|((~II32659));
assign g21356 = (g9488&g20355);
assign g30828 = ((~II40736));
assign g28439 = (g28128&g9242);
assign II13186 = ((~g1088));
assign g23245 = ((~II30188));
assign gbuf124 = (g1657);
assign g13969 = (g7652&g12891);
assign g16672 = ((~g15962)&(~g14703)&(~g15923));
assign II25597 = ((~g18074))|((~II25595));
assign g13738 = (g6887&g12545);
assign g29556 = ((~II38940));
assign g24267 = ((~II31475));
assign g4948 = ((~g1754));
assign II40107 = ((~g30343));
assign g19369 = ((~II25778));
assign g7053 = ((~II14891));
assign g22092 = ((~g21354)&(~g19639));
assign g27408 = ((~g27012))|((~g5473));
assign g19351 = (g16924&g16599&g14301);
assign II35109 = ((~g26676));
assign g12376 = (g7974&g8949);
assign gbuf92 = (g1059);
assign II31426 = ((~g22615));
assign g19648 = (g2072&g18814);
assign g23867 = ((~II31121));
assign g19175 = ((~II25386));
assign g26640 = ((~g25787));
assign g12442 = ((~II19602));
assign g10512 = (g7162&g5061);
assign g28078 = ((~II36679));
assign g20779 = ((~g20255))|((~g3722));
assign g10675 = (g7488&g5323);
assign II29478 = ((~g21006));
assign g19874 = (g1372&g18930);
assign g28359 = ((~II37252));
assign g18936 = ((~g15635));
assign II19784 = ((~g8726));
assign II35407 = ((~g27145));
assign g28834 = (g5751&g28483);
assign g16439 = ((~g13082))|((~g2912));
assign g10294 = (g3410&g4629);
assign g15178 = (g640&g12651);
assign g17161 = (g7712&g14183);
assign g29628 = ((~II39002));
assign g9100 = (g7265&g7697);
assign g3616 = ((~II13203));
assign g4035 = ((~g845));
assign g29791 = ((~g29490)&(~g29243));
assign g12078 = ((~g11422));
assign g5804 = ((~g237));
assign II24678 = ((~g6305))|((~II24677));
assign g5787 = (g1712&g1747);
assign g7161 = ((~II14917));
assign g10639 = (g7303&g5275);
assign g21639 = (g3398&g20500);
assign g9894 = (g6448&g4112);
assign II33539 = ((~g24458));
assign g19699 = (g660&g18840);
assign g27913 = (g4017&g27401);
assign g13134 = ((~g9676))|((~g6980));
assign II15549 = ((~g6574));
assign g22885 = ((~g21863))|((~g21859))|((~g21885));
assign g20996 = ((~g19810)&(~g15486));
assign II16185 = ((~g5415));
assign g27582 = ((~g26944)&(~g24731));
assign g26282 = ((~II34244));
assign g19704 = (g4243&g17520);
assign g19972 = ((~II26420));
assign II15359 = ((~g2858));
assign g28007 = ((~II36502));
assign II16785 = ((~g7053));
assign g23310 = ((~II30383));
assign II24554 = ((~g6163))|((~II24553));
assign g24243 = ((~g17097)&(~g22333));
assign g22588 = ((~g21099));
assign II31841 = ((~g23607));
assign g30019 = ((~g29538)&(~g29952));
assign g27002 = (g23335&g26571);
assign g28552 = ((~II37481));
assign g4662 = ((~g1400));
assign II37228 = ((~g28194));
assign g29283 = ((~g28799));
assign g11707 = ((~g9534))|((~g3366));
assign g12108 = ((~g10314)&(~g10392)&(~g10454));
assign g28859 = ((~g28413));
assign g11762 = ((~g10915));
assign II37973 = ((~g28556));
assign g28069 = ((~II36650));
assign II31562 = ((~g23594));
assign g18898 = ((~g15483));
assign g5170 = ((~g1772));
assign g27271 = ((~g26999)&(~g26299));
assign g10825 = ((~II17670));
assign g26450 = (g5204&g25805);
assign g19560 = (g8065&g17259);
assign g16829 = ((~g14956)&(~g12564));
assign g15546 = (g5057&g13238);
assign g14234 = ((~g12008));
assign g19476 = (g16913&g14849&g14811);
assign g11069 = ((~g8257));
assign II38342 = ((~g28886));
assign II33532 = ((~g24507));
assign g9873 = ((~II16867));
assign g13243 = ((~g9965));
assign g21819 = (g20184)|(g20148)|(g18629)|(g19109);
assign g25933 = ((~g24989))|((~g5512));
assign g8577 = ((~g3866))|((~g3834));
assign g24897 = ((~II32625))|((~II32626));
assign g8065 = ((~g831));
assign g19884 = (g2734&g18938);
assign II23791 = ((~g15951));
assign g6227 = ((~g3100));
assign g24310 = ((~II31604));
assign g30030 = ((~g24676)&(~g29923));
assign gbuf43 = (g372);
assign II29610 = ((~g21052));
assign g21946 = ((~II28464));
assign II23880 = ((~g9187))|((~II23878));
assign g19096 = ((~g18980));
assign II13228 = ((~g2476));
assign g8526 = (g6574&g1648);
assign II32704 = ((~g23357));
assign g13065 = ((~g9822))|((~g7358));
assign g25983 = ((~II33801));
assign II33689 = ((~g25074));
assign g25827 = ((~II33667));
assign g20436 = ((~g17704));
assign g19277 = ((~II25579))|((~II25580));
assign g9925 = (g3566&g4165);
assign II27328 = ((~g19369));
assign g10870 = ((~II17727));
assign g25419 = ((~g24812));
assign g5763 = ((~g912));
assign II35497 = ((~g27158));
assign II22667 = ((~g14642));
assign II40110 = ((~g30357));
assign II21982 = ((~g13137));
assign g5041 = ((~g1078));
assign g24581 = ((~II32137));
assign g11059 = ((~II17978));
assign II31133 = ((~g22185));
assign II19891 = ((~g10708));
assign g8877 = ((~II16141));
assign g25699 = ((~g24613)&(~g24506));
assign g10018 = ((~II16990));
assign g27228 = ((~II35521));
assign g15363 = ((~II21632));
assign g13368 = (g5795&g11404);
assign g10415 = (g7426&g4879);
assign g6000 = ((~II14472));
assign g20366 = ((~g17451));
assign g29703 = ((~g29583)&(~g1917));
assign II24560 = ((~g13611));
assign g4564 = ((~g2237));
assign g25010 = ((~g23694))|((~g6713));
assign II34111 = ((~g25223));
assign gbuf193 = (g2462);
assign II40724 = ((~g30656));
assign II21429 = ((~g13027));
assign g19270 = ((~II25557));
assign g26958 = (g6184&g26538);
assign II18488 = ((~g8840));
assign g25086 = (g23444&g10880);
assign g11216 = ((~II18142));
assign g13123 = ((~g9534))|((~g6678));
assign II16172 = ((~g5413));
assign g7423 = ((~g2533));
assign g29270 = ((~II38391));
assign g12904 = ((~II19961));
assign g10036 = (g6912&g4228);
assign g21180 = (g20150&g14565);
assign g30724 = ((~II40462));
assign g27973 = ((~II36444));
assign II18527 = ((~g10017));
assign g9228 = ((~g7667));
assign g13033 = ((~g10797));
assign g28656 = ((~g27772)&(~g27358));
assign II37716 = ((~g28540));
assign g22645 = ((~g21125));
assign II21609 = ((~g11692));
assign g13835 = (g7461&g12600);
assign g11785 = ((~g9464)&(~g9583)&(~g9663));
assign g13701 = (g6623&g12536);
assign g10147 = ((~g7788))|((~g3522));
assign g28281 = ((~II37092));
assign II38278 = ((~g28963));
assign g20425 = ((~g17664));
assign g22875 = ((~g21884));
assign g9722 = (g3566&g3966);
assign g24938 = (g24084&g18967);
assign g10378 = (g6751&g4783);
assign g27729 = (g27435&g19322);
assign g6099 = ((~II14612));
assign g18788 = ((~g15052));
assign II15779 = ((~g6000));
assign g8382 = ((~II15584));
assign g11537 = ((~II18587));
assign g30392 = (g30237&g8968);
assign II19855 = ((~g10723));
assign g24859 = ((~g16390)&(~g24253));
assign g24378 = ((~II31808));
assign g29736 = ((~g29583)&(~g25444));
assign g28123 = (g27622&g10337);
assign g9355 = ((~g7639));
assign II24308 = ((~g15274))|((~II24306));
assign g22754 = (g14342&g21612);
assign g16008 = (g5504&g11735);
assign g19851 = (g2040&g18919);
assign g18649 = (g14776&g14837&g13657&g16189);
assign g9027 = ((~g5679));
assign g17258 = ((~g16053));
assign II21329 = ((~g11766));
assign II40245 = ((~g30381));
assign g24386 = ((~II31832));
assign II31205 = ((~g22002));
assign g21599 = ((~II28130));
assign II27565 = ((~g19987));
assign g28678 = ((~II37581));
assign g20920 = ((~g19691)&(~g19726));
assign II38920 = ((~g29204));
assign g28349 = ((~g15595)&(~g28051));
assign g27820 = ((~II36283));
assign g26708 = ((~II34731));
assign g12932 = ((~g8968));
assign g20185 = (g16313&g13797&II26624);
assign g7795 = ((~g2992)&(~g2991));
assign g11501 = ((~II18479));
assign g11573 = ((~II18695));
assign g30058 = ((~g29968)&(~g13395));
assign g19238 = ((~II25489));
assign II38088 = ((~g28361));
assign g24208 = ((~g16969)&(~g22235));
assign g15711 = ((~II21959));
assign g26815 = ((~g15350)&(~g26311));
assign g28581 = ((~g27817));
assign g12531 = (g7868&g9146);
assign g24371 = ((~II31787));
assign II16472 = ((~g7901));
assign g29965 = (g29756&g11961);
assign g13052 = ((~g9822))|((~g7230));
assign g26869 = ((~g26458)&(~g5642));
assign g15757 = ((~g11622))|((~g12392));
assign g29143 = ((~II38172));
assign g30361 = (g30203&g8440);
assign g23301 = ((~II30356));
assign g25289 = (g5631&g24834);
assign g26566 = ((~g25540));
assign g22650 = (g14033&g21518);
assign g8018 = ((~g2969));
assign g5982 = ((~g785));
assign g8944 = ((~II16244));
assign g24782 = ((~g16160)&(~g24221));
assign II33498 = ((~g25036));
assign II35058 = ((~g26137))|((~II35057));
assign g8909 = ((~II16193));
assign II38172 = ((~g29085));
assign g24841 = (g12974&g24177);
assign II34579 = ((~g25452));
assign II35373 = ((~g26189));
assign g20901 = ((~g19660)&(~g17508));
assign g14895 = ((~g12193));
assign g12691 = ((~g8805));
assign g29936 = ((~g16049)&(~g29790));
assign g24223 = ((~g17018)&(~g22273));
assign g17486 = (g4091&g16014);
assign g20644 = ((~II27235));
assign II18740 = ((~g8978));
assign II35035 = ((~g26087))|((~II35034));
assign g5552 = ((~II14034));
assign g27414 = ((~g26770)&(~g25187));
assign g18991 = ((~II25061));
assign II24500 = ((~g6626))|((~g14044));
assign g16198 = (g5762&g11866);
assign g26609 = ((~g25672));
assign g26173 = ((~II34071));
assign g21012 = ((~II27565));
assign II38668 = ((~g29168));
assign II31937 = ((~g24079));
assign g11956 = ((~g10078)&(~g10169)&(~g10256));
assign g22363 = (g776&g21199);
assign II37729 = ((~g28567));
assign II24123 = ((~g6290))|((~g14201));
assign g21106 = ((~g20053)&(~g20090)&(~g20112));
assign g5949 = (g2412&g2399);
assign g14794 = ((~g11848));
assign II20586 = ((~g11606));
assign g13460 = ((~II20679));
assign II28201 = ((~g20025));
assign g5668 = ((~g299));
assign g7528 = ((~g3151)&(~g3142)&(~g3147));
assign II35003 = ((~g26592));
assign g25147 = ((~II32919));
assign g14298 = ((~II21149));
assign II36598 = ((~g27294));
assign II36499 = ((~g27268));
assign g25123 = ((~II32857));
assign g8856 = ((~II16104));
assign g23182 = ((~II29999));
assign g13486 = (g6023&g12212);
assign g24475 = ((~g24014))|((~g3806));
assign II30011 = ((~g22758));
assign II33399 = ((~g25018));
assign g15354 = ((~g12259));
assign II15836 = ((~g3366));
assign II40919 = ((~g30781));
assign g26019 = ((~II33909));
assign II27146 = ((~g19838));
assign g12708 = ((~II19800));
assign II30161 = ((~g22133));
assign g6230 = ((~II14709));
assign g29347 = ((~g28340)&(~g28729));
assign g25124 = ((~II32860));
assign g25215 = ((~g24755)&(~g23564));
assign g12186 = (g8093&g8805);
assign g29421 = ((~II38644));
assign g27540 = ((~II35926));
assign g24778 = ((~II32309))|((~II32310));
assign g27288 = ((~g27022)&(~g26343));
assign g16494 = ((~II22584));
assign g10269 = (g3834&g4578);
assign g17050 = ((~II23035))|((~II23036));
assign g22841 = (g7583&g21902);
assign g10260 = (g3774&g2489);
assign g29563 = ((~II38951));
assign g17785 = ((~II23860));
assign g22774 = ((~II29536));
assign g15635 = ((~II21888));
assign g25388 = (g5971&g24630);
assign II18799 = ((~g11410))|((~g11331));
assign g25029 = ((~g23923))|((~g6486));
assign g17531 = ((~II23619));
assign g29685 = ((~g29564)&(~g29341));
assign g21234 = (g19608&g14849&g16686);
assign g25688 = ((~II33514));
assign g23129 = (g21823)|(g21820);
assign g21362 = (g15096&g20363);
assign II27942 = ((~g19157));
assign II35083 = ((~g26665));
assign g21074 = ((~g19929)&(~g18245));
assign g27200 = ((~II35437));
assign g10470 = (g3774&g2510);
assign g17148 = ((~II23172))|((~II23173));
assign g15718 = ((~g13286))|((~g12354));
assign g10661 = (g7195&g1997);
assign g26477 = (g5269&g25841);
assign II15833 = ((~g3338));
assign g8197 = ((~g154));
assign g5706 = ((~g231));
assign g24431 = (g17124&g24153&g13637);
assign II39164 = ((~g29621));
assign II40715 = ((~g30653));
assign g28923 = (g28625&g9338);
assign g22192 = ((~g21521)&(~g19856));
assign g24053 = ((~II31270));
assign II29435 = ((~g20992));
assign g24406 = ((~II31892));
assign II23760 = ((~g15897));
assign g10258 = (g6838&g4567);
assign g8485 = (g3254&g255);
assign II29007 = ((~g21760));
assign II37659 = ((~g28437));
assign g7576 = ((~g468));
assign g26232 = ((~II34172));
assign g10319 = (g3678&g4693);
assign g20780 = ((~II27369));
assign g8467 = (g6519&g930);
assign II40916 = ((~g30777));
assign g30974 = ((~II41096));
assign g27455 = ((~g23127)&(~g26758)&(~g24431));
assign II14413 = ((~g3233));
assign II27358 = ((~g19369));
assign g7878 = ((~g3056));
assign g19045 = ((~II25198));
assign g27207 = ((~II35458));
assign g26658 = ((~g25865));
assign g7549 = ((~g3028));
assign g20455 = ((~g17791));
assign g20345 = ((~g17387));
assign II40651 = ((~g30574));
assign g21903 = ((~g20008))|((~g3013));
assign g28661 = ((~g27775)&(~g27371));
assign g16359 = (g5909&g11996);
assign g11864 = ((~g9778)&(~g9906)&(~g10042));
assign g13127 = ((~g9822))|((~g7230));
assign g14222 = ((~g12933));
assign g20285 = (g16846&g8103);
assign g16024 = ((~g12702));
assign g28192 = ((~g27372)&(~g26866));
assign g21122 = (g20140&g12279);
assign II29142 = ((~g20682));
assign II26916 = ((~g17271));
assign II20848 = ((~g13194));
assign g23408 = ((~g22606)&(~g21494));
assign II37946 = ((~g28529));
assign II26383 = (g18483&g18405&g18331);
assign g25664 = ((~II33488));
assign g13026 = ((~g9534))|((~g6678));
assign g28073 = (g27595&g10109);
assign g10754 = ((~g4848));
assign g17351 = ((~g16152));
assign g11736 = ((~g10862));
assign II14478 = ((~g3213));
assign g19759 = (g2707&g18863);
assign g29316 = ((~II38477));
assign g27661 = (g26841&g11173);
assign g30478 = (g30187&g11344);
assign g5227 = ((~g2805));
assign II37296 = ((~g27827))|((~II37295));
assign g24367 = ((~II31775));
assign II33402 = ((~g24448));
assign g21850 = ((~g17979))|((~g19187))|((~g19191));
assign g19795 = (g2707&g18880);
assign g25681 = ((~II33507));
assign g27071 = (g23353&g26632);
assign II23152 = ((~g9427))|((~g14061));
assign II22981 = ((~g15274))|((~g14106));
assign g19940 = (g2753&g18973);
assign g8488 = (g3410&g933);
assign g30326 = ((~II39821));
assign II20562 = ((~g11786));
assign II19852 = ((~g10679));
assign g12438 = ((~g10846));
assign g18368 = ((~g14286));
assign g5776 = ((~g1597));
assign g26165 = ((~II34059));
assign g28237 = ((~II36960));
assign II37814 = ((~g28388))|((~II37813));
assign II25880 = ((~g776))|((~g17914));
assign g14182 = (g7733&g12969);
assign g15263 = ((~g12369));
assign g26726 = ((~II34785));
assign II36516 = ((~g27273));
assign g24763 = ((~II32281));
assign g10949 = ((~II17846));
assign g9623 = ((~II16720));
assign g28025 = ((~II36542));
assign g16358 = (g5908&g11995);
assign g6032 = ((~g897));
assign II29301 = ((~g20944));
assign g15890 = ((~g11600));
assign g28477 = (g18341&g28174);
assign g8141 = ((~g834));
assign II33646 = ((~g24468));
assign II18206 = ((~g4202))|((~II18204));
assign g27303 = ((~g27043)&(~g26380));
assign g15174 = ((~g12136));
assign g26037 = ((~g25311)&(~g18407));
assign g15296 = ((~g11882));
assign II40212 = ((~g30471));
assign II25234 = ((~g16906));
assign g11199 = ((~II18121));
assign g4549 = ((~g2081));
assign g27196 = ((~II35425));
assign g12876 = (II19937&II19938);
assign II38205 = ((~g28924));
assign g21965 = ((~II28521));
assign II35727 = ((~g26902));
assign g10813 = ((~II17658));
assign II29533 = ((~g21026));
assign g17717 = (g4587&g15385);
assign g10154 = (g3566&g4401);
assign II38524 = ((~g28788));
assign II31745 = ((~g23669));
assign g26120 = ((~g23694))|((~g25369));
assign g30105 = (g29861&g11364);
assign g9903 = (g6678&g4121);
assign II28119 = ((~g19957));
assign g26644 = ((~g25805));
assign g16460 = (g5998&g12175);
assign g27266 = ((~g26994)&(~g26289));
assign g26239 = ((~II34183));
assign II29317 = ((~g20949));
assign g16389 = (g5936&g12040);
assign g10316 = ((~II17278));
assign g12815 = ((~g8856));
assign g24921 = (g24073&g18951);
assign II31282 = ((~g22263));
assign g25227 = ((~g24775)&(~g23586));
assign g23170 = ((~II29963));
assign g8518 = (g3254&g273);
assign g27937 = ((~g16321)&(~g27666));
assign g24522 = ((~g15476)&(~g23860));
assign II37113 = ((~g28044));
assign II21809 = ((~g13125));
assign II40955 = ((~g30734));
assign g27281 = ((~g27009)&(~g26326));
assign g22077 = ((~g21341)&(~g19620));
assign g27683 = ((~II36060));
assign g28110 = ((~II36761));
assign g28680 = ((~II37587));
assign g27802 = ((~g6087)&(~g27632)&(~g25330));
assign g30460 = (g30155&g11231);
assign g25589 = ((~g20850)&(~g24433));
assign II24992 = ((~g14936));
assign g14863 = ((~g12169));
assign g28413 = ((~g24695)&(~g27809));
assign g26158 = (g679&g25937);
assign g9174 = ((~g5932));
assign II25489 = ((~g18906));
assign g21870 = ((~g18497))|((~g19223))|((~g19231));
assign g26855 = ((~II35014));
assign gbuf164 = (g1929);
assign g21261 = (g19641)|(g16770)|(g14863);
assign g5675 = ((~g302));
assign g5058 = ((~g1402));
assign g11796 = ((~g10980));
assign II23144 = ((~g13991))|((~II23142));
assign g27105 = (g22134&g26656);
assign g18909 = ((~g15528));
assign gbuf188 = (g2440);
assign II30359 = ((~g22934));
assign g11256 = ((~II18184));
assign g27419 = ((~II35759));
assign g21665 = ((~g20507)&(~g18352));
assign g12112 = ((~g10321)&(~g10397)&(~g10460));
assign g26860 = (g5774&g26070);
assign g24342 = ((~II31700));
assign II32686 = ((~g18155))|((~g24028));
assign g14957 = (g4015&g13152);
assign II39936 = ((~g30299));
assign g20927 = ((~g19710)&(~g17600));
assign g11190 = ((~g3999));
assign II30769 = ((~g22078));
assign II18019 = ((~g6945));
assign g13303 = ((~g10263));
assign g11998 = ((~g11312));
assign II36755 = ((~g27336));
assign II32847 = ((~g24083));
assign g15314 = ((~II21583));
assign g11933 = ((~g11210));
assign g25053 = ((~g23923))|((~g6486));
assign g18968 = ((~g13904)&(~g12330));
assign g25194 = ((~g24514)&(~g10238));
assign g29118 = ((~II38122));
assign g11297 = ((~II18247));
assign II24696 = ((~g14374))|((~II24694));
assign II35334 = ((~g26106));
assign g21618 = ((~g20016)&(~g14079)&(~g14165));
assign II25355 = ((~g18669));
assign g27345 = ((~g27101)&(~g26479));
assign g10843 = ((~II17692));
assign g29771 = ((~g29472)&(~g29200));
assign g5012 = ((~g2786));
assign g28839 = ((~II37808));
assign g8563 = ((~g3710))|((~g3678));
assign II25782 = ((~g1444))|((~II25781));
assign g5256 = ((~g1994));
assign g27980 = ((~g16428)&(~g27681));
assign g25738 = ((~II33567));
assign g29565 = (g28795&g29394);
assign g6189 = ((~g1934));
assign g21894 = ((~g19317)&(~g19356));
assign g30563 = ((~II40269));
assign g27075 = ((~II35254));
assign g23068 = ((~II29817));
assign g30887 = ((~II40913));
assign g10792 = ((~II17637));
assign II36630 = ((~g27303));
assign g25062 = ((~g24014))|((~g7303));
assign g27535 = ((~II35919));
assign g24182 = ((~g16953)&(~g22223));
assign II37740 = ((~g28595));
assign g22727 = (g14238&g21590);
assign g30525 = ((~II40155));
assign g28687 = ((~II37608));
assign g25075 = ((~g13880)&(~g23483));
assign g4406 = ((~g1809));
assign g17737 = (g4626&g15404);
assign g21222 = ((~II27785));
assign g14205 = ((~g11992));
assign g8400 = ((~II15602));
assign g13204 = ((~g9626));
assign g16188 = (g5755&g11858);
assign II15915 = ((~g3878));
assign g25072 = ((~g24014))|((~g7303));
assign g8212 = ((~g837));
assign g21411 = (g9649&g20403);
assign II30748 = ((~g21969));
assign g13148 = ((~g9170));
assign g22796 = ((~II29572));
assign g18458 = ((~II24486))|((~II24487));
assign g30119 = ((~II39622));
assign g21152 = (g19357&g19334&II27711);
assign II27488 = ((~g20310));
assign g5407 = ((~II13937));
assign II23172 = ((~g9471))|((~II23171));
assign g28498 = ((~II37459));
assign g13346 = ((~II20425));
assign g14752 = (g7891&g13130);
assign II26796 = ((~g17224));
assign g12852 = ((~g8439)&(~g8467)&(~g8488));
assign g29776 = ((~g29477)&(~g29220));
assign g19978 = ((~II26426));
assign II41065 = ((~g30927))|((~II41064));
assign g16546 = ((~g14366));
assign g10106 = (g6448&g432);
assign II21304 = ((~g11927));
assign II39368 = ((~g29767))|((~II39367));
assign g28259 = ((~II37026));
assign g28607 = ((~II37508));
assign g11411 = ((~II18375));
assign g24804 = (g12945&g24152);
assign g20968 = ((~g19767)&(~g17736));
assign g5745 = ((~g2200));
assign g12051 = ((~g11376));
assign g20433 = ((~g17691));
assign II30362 = ((~g22636));
assign II19240 = ((~g9341));
assign g17850 = ((~II23911));
assign II25890 = ((~g18453))|((~II25888));
assign g17150 = ((~II23180))|((~II23181));
assign g29756 = ((~g16284)&(~g29614));
assign g23049 = ((~g21590));
assign g20919 = ((~g19688)&(~g17555));
assign g13273 = ((~g10130));
assign II32583 = ((~g23330));
assign g29666 = ((~g29577));
assign g27024 = (g23372&g26593);
assign g8631 = (g6751&g6974);
assign II30813 = ((~g22091));
assign g9038 = ((~II16357));
assign g11800 = ((~g9523)&(~g9634)&(~g9762));
assign g21490 = (g15296&g20453);
assign g27706 = ((~II36129));
assign g19191 = (g17807)|(g17887);
assign g24147 = ((~g22512));
assign g17128 = (g7479&g15678);
assign g24444 = ((~g23694))|((~g3462));
assign g20539 = ((~II26980));
assign g14776 = ((~g12033));
assign g12506 = ((~g8287))|((~g6713));
assign g28212 = ((~II36885));
assign g5637 = ((~II14091));
assign g21983 = ((~g19255))|((~g21139))|((~g19294));
assign g11971 = ((~g11274));
assign g29704 = ((~II39164));
assign g9062 = (g5438&g7626);
assign g29164 = ((~II38235));
assign g22143 = ((~g21403)&(~g19729));
assign II38591 = ((~g28987));
assign II39625 = ((~g30076));
assign g25796 = ((~II33633));
assign g20084 = (g17969&g3158);
assign II29459 = ((~g21000));
assign g17223 = ((~g15981)&(~g14737));
assign g18827 = ((~g15204));
assign g24413 = ((~II31913));
assign II34716 = ((~g26215));
assign g30253 = ((~g16222)&(~g30087));
assign II29582 = ((~g21044));
assign g26783 = (g26073&g19326);
assign II17645 = ((~g6288));
assign g19623 = (g4000&g17384);
assign g24233 = ((~II31417));
assign II35737 = ((~g26915));
assign g30890 = ((~II40922));
assign II24325 = ((~g14124))|((~g9857));
assign g12611 = ((~II19759));
assign g22183 = ((~g21488)&(~g19822));
assign g16382 = (g5927&g12022);
assign g18897 = ((~g15480));
assign g21497 = (g3006&g20456);
assign II38330 = ((~g29120));
assign g5880 = ((~g2180));
assign g23610 = (g4085&g22506);
assign g14011 = ((~g11896));
assign g20586 = ((~II27083));
assign II34827 = ((~g26315));
assign g7841 = ((~g630));
assign g29426 = ((~II38659));
assign g16583 = ((~g14507)&(~g14601));
assign g19912 = (g2753&g18955);
assign II30047 = ((~g22107));
assign g8276 = ((~g3253));
assign g18415 = ((~g15783));
assign g13001 = ((~g8553)&(~g8562)&(~g8570));
assign g27604 = ((~g27157));
assign g11855 = ((~g9761)&(~g9889)&(~g10009));
assign II30386 = ((~g22839));
assign g15578 = ((~g12346));
assign g11599 = ((~II18773));
assign g22250 = (g21752&g12225);
assign g4845 = ((~g2112));
assign g11979 = ((~g10114)&(~g10202)&(~g10288));
assign g29353 = ((~g29126)&(~g17001));
assign g9199 = ((~II16479));
assign g27504 = ((~g26918)&(~g24656));
assign g9920 = (g6980&g4150);
assign II22715 = ((~g14711));
assign g13456 = ((~II20667));
assign g23524 = ((~II30568));
assign g10061 = (g6574&g4272);
assign g9081 = (g7015&g7661);
assign II19648 = ((~g10855));
assign g13503 = (g6037&g12265);
assign II35488 = ((~g26819));
assign g26222 = ((~II34156));
assign gbuf84 = (g975);
assign II16071 = ((~g5395));
assign II16068 = ((~g5438));
assign g10525 = (g3678&g5098);
assign II30143 = ((~g22678));
assign g11048 = ((~II17963));
assign g26814 = ((~g15338)&(~g26303));
assign II39361 = ((~g15880))|((~II39359));
assign II38059 = ((~g28352));
assign II23218 = ((~g9613))|((~II23217));
assign g30899 = ((~II40949));
assign g28982 = ((~g28665)&(~g28670));
assign g8924 = ((~II16212));
assign II28727 = ((~g21887))|((~II28726));
assign g30810 = ((~II40682));
assign II39815 = ((~g30313));
assign g19592 = (g8236&g17333);
assign II23911 = ((~g14985));
assign g23012 = ((~g21505));
assign g15701 = ((~II21949));
assign g30512 = ((~II40116));
assign g24276 = ((~II31502));
assign II16031 = ((~g3878));
assign g28199 = ((~g27250)&(~g10024));
assign II31640 = ((~g23691));
assign g14378 = ((~g12100));
assign g7916 = ((~g2935));
assign II32595 = ((~g18014))|((~g23938));
assign g25158 = ((~II32952));
assign g21219 = ((~g19253)&(~g19243));
assign II34785 = ((~g26448));
assign g22546 = (g13886&g21404);
assign II39270 = ((~g29700));
assign g21491 = ((~II28027));
assign g13864 = ((~g11767));
assign g13290 = ((~II20347));
assign g7140 = ((~g2170));
assign g20379 = ((~g17490));
assign II33511 = ((~g24456));
assign g27595 = ((~g27149));
assign g30004 = (g29926&g22295);
assign II38211 = ((~g29095));
assign II34803 = ((~g26248));
assign II31667 = ((~g23452));
assign g19390 = ((~II25816));
assign g8260 = ((~II15448));
assign II32365 = ((~g24009));
assign II25412 = ((~g18820));
assign g18578 = ((~II24668))|((~II24669));
assign II16499 = ((~g7901));
assign g9450 = ((~II16633));
assign g15065 = ((~g12291));
assign g7141 = ((~g2195));
assign g27246 = (g26988&g16676);
assign II26874 = ((~g17236));
assign g15880 = ((~g11624));
assign g8997 = ((~II16315));
assign g27191 = ((~II35410));
assign II17311 = ((~g3900));
assign II34405 = ((~g25933));
assign g26790 = (g26079&g19353);
assign g22445 = ((~II28991));
assign II28470 = ((~g20984));
assign g12533 = ((~g8673));
assign II13113 = ((~g11));
assign g26691 = ((~II34680));
assign II35141 = ((~g26666));
assign g11008 = ((~II17919));
assign g26055 = ((~g25881)&(~g24974));
assign II23256 = ((~g9795))|((~g14205));
assign II40799 = ((~g30723));
assign II26895 = ((~g17247));
assign g23770 = (g22921&g20454);
assign g14975 = (g4047&g13154);
assign g22559 = ((~II29119));
assign II18091 = ((~g7195));
assign g7661 = ((~g1694));
assign g22591 = ((~II29165));
assign g29807 = ((~II39273));
assign g11543 = ((~II18605));
assign g28434 = (g26114&g28159);
assign g23911 = ((~II31181));
assign II22657 = ((~g14657));
assign II30704 = ((~g22058));
assign g30915 = ((~II40997));
assign g13111 = ((~g8601)&(~g8612)&(~g8621));
assign g7877 = ((~g3046));
assign g6084 = ((~II14599));
assign II18199 = ((~g7876))|((~II18197));
assign II25195 = ((~g18932));
assign g29234 = (g9427&g28804);
assign g23738 = ((~II30928));
assign II25406 = ((~g18804));
assign g19562 = (g8076&g17265);
assign II19510 = ((~g10574));
assign II40054 = ((~g30258));
assign II18114 = ((~g3997))|((~II18113));
assign g21321 = (g9248&g20317);
assign g16804 = ((~g15803));
assign g11611 = ((~II18787));
assign g25360 = (g24664&g18200);
assign g10386 = (g6980&g4803);
assign g22512 = ((~II29058));
assign II27416 = ((~g19420));
assign g11827 = ((~g11032));
assign II30632 = ((~g22035));
assign g12346 = ((~II19513));
assign II16796 = ((~g5556));
assign g20392 = ((~g17545));
assign II36147 = ((~g27560));
assign g25510 = ((~II33338));
assign II33445 = ((~g25026));
assign g21343 = (g9161&g20344);
assign g30897 = ((~II40943));
assign II22705 = ((~g13348))|((~g15661));
assign g21056 = ((~g19905)&(~g18130));
assign g5695 = ((~II14143));
assign II30173 = ((~g22656));
assign II20062 = ((~g10480));
assign g28935 = (g14177&g28646);
assign II17771 = ((~g8107));
assign g26316 = (g4717&g25562);
assign g23074 = ((~g21623));
assign g5260 = ((~g2104));
assign g16309 = (g1205&g11945);
assign g22176 = ((~II28712));
assign g18906 = ((~g13855)&(~g12186));
assign II37152 = ((~g28109));
assign II31574 = ((~g23736));
assign g12324 = ((~g10626)&(~g10661)&(~g10681));
assign II31529 = ((~g23729));
assign g20625 = ((~II27200));
assign g17511 = ((~II23599));
assign g30337 = (g30199&g8354);
assign II36591 = ((~g27529))|((~g14885));
assign g19326 = ((~g16640));
assign g29130 = (g28397&g22221);
assign g22065 = ((~g21330)&(~g19599));
assign g24305 = ((~II31589));
assign g3248 = ((~II13140));
assign g10592 = (g7391&g5210);
assign g11695 = ((~g9968))|((~g3834));
assign g17749 = ((~II23824));
assign g28099 = ((~II36728));
assign g28230 = ((~II36939));
assign g18290 = ((~II24291))|((~II24292));
assign II18695 = ((~g11054));
assign II39333 = ((~g29751))|((~II39331));
assign g19617 = (g3969&g17366);
assign g24112 = ((~g22445));
assign g20477 = ((~g17962));
assign g5822 = ((~g1606));
assign II30654 = ((~g22042));
assign g23570 = ((~II30642));
assign g22560 = ((~II29122));
assign g16846 = ((~g15903));
assign g11361 = ((~II18317));
assign g30448 = (g30151&g11148);
assign g7591 = ((~g1496));
assign g30823 = ((~II40721));
assign g20117 = (g16189&g13706&II26561);
assign g16472 = ((~II22518));
assign II39121 = ((~g29579));
assign g12752 = ((~II19816));
assign g28023 = ((~II36536));
assign g25339 = ((~g24887));
assign II30395 = ((~g22253));
assign g30859 = ((~II40829));
assign g30279 = ((~g16424)&(~g30113));
assign II27402 = ((~g19420));
assign g16323 = (g5878&g11959);
assign g26068 = (g2138&g25324);
assign g14884 = (g8169&g12548);
assign g25183 = (g24958)|(g24893);
assign II37167 = ((~g28121));
assign g11453 = ((~II18417));
assign II23421 = ((~g15791));
assign g7809 = ((~g1702));
assign g9765 = (g5438&g417);
assign g19674 = (g2020&g18830);
assign g27143 = ((~g26150));
assign II35817 = ((~g26922));
assign g12998 = ((~g9044));
assign g25383 = ((~g24766));
assign g5757 = (g337&g383);
assign II25985 = ((~g16718));
assign g5375 = ((~g2812));
assign g22739 = ((~g16164))|((~g21285));
assign g21805 = (g16679&g19578&g14776);
assign g15506 = (g4845&g12833);
assign g30008 = (g29919&g22334);
assign g25036 = ((~g23748))|((~g7015));
assign g24812 = ((~II32379))|((~II32380));
assign g10626 = (g7053&g1994);
assign g7079 = ((~g2040));
assign II36954 = ((~g28010));
assign II26990 = ((~g19145));
assign g24179 = ((~g16923)&(~g22214));
assign II20791 = ((~g13149));
assign II15955 = ((~g3878));
assign g10746 = ((~g3866))|((~g7426));
assign g22123 = ((~g21379)&(~g19693));
assign g22934 = ((~II29715));
assign II39859 = ((~g30277));
assign II36779 = ((~g27577))|((~g15151));
assign g6184 = ((~g1372));
assign II30077 = ((~g22675));
assign g19384 = ((~g17132));
assign g24165 = ((~g22567));
assign g16619 = ((~g14601));
assign II33864 = ((~g25796));
assign g8559 = (g3410&g897);
assign g27687 = ((~II36072));
assign g13324 = ((~g10316));
assign g26264 = ((~II34220));
assign II27900 = ((~g19096));
assign g17969 = ((~g15841));
assign g18975 = ((~g13944)&(~g12353));
assign II19523 = ((~g10500));
assign g19079 = (g14797&g18692&g16142&g16189);
assign g4228 = ((~g706));
assign g27256 = ((~g26970)&(~g26234));
assign g19695 = (g4214&g17496);
assign g30956 = ((~g30919)&(~g30946));
assign II30869 = ((~g22881))|((~II30868));
assign g5279 = ((~g2679));
assign II27143 = ((~g19763));
assign g27558 = ((~g24993)&(~g24691)&(~g26791));
assign g19758 = (g2714&g18862);
assign g8542 = (g6838&g2261);
assign g22635 = ((~II29235));
assign g19381 = (g16924&g16578&g14395);
assign g22364 = ((~g21189));
assign g29045 = ((~g9232))|((~g28512));
assign g30249 = ((~g16158)&(~g30082));
assign g16230 = ((~g10952)&(~g6220)&(~g12539));
assign g30262 = ((~g16343)&(~g30096));
assign g20619 = ((~II27182));
assign g29544 = ((~II38920));
assign g25332 = ((~g24900));
assign II28093 = ((~g19957));
assign g18523 = ((~II24582));
assign g22764 = (g18374&g21623);
assign g12282 = ((~II19452));
assign g26457 = (g5213&g25814);
assign g19155 = (g17200&g8614);
assign g8074 = ((~g1172));
assign g7769 = ((~g323));
assign g12419 = (g8028&g9006);
assign g10808 = ((~II17653));
assign g10079 = (g3722&g4304);
assign g30544 = ((~II40212));
assign g11916 = ((~g9954)&(~g10077)&(~g10168));
assign g21640 = ((~II28169));
assign II40629 = ((~g30594))|((~II40627));
assign g29496 = ((~II38804));
assign g22131 = ((~g21394)&(~g19712));
assign g13564 = ((~g12711))|((~g3722));
assign II16276 = ((~g5512));
assign g23196 = ((~II30041));
assign g4354 = ((~g711));
assign g24356 = ((~II31742));
assign g25135 = ((~II32883));
assign g26107 = ((~g6068)&(~g24183)&(~g25383));
assign g30269 = ((~g16386)&(~g30103));
assign g22236 = ((~g20641));
assign g28720 = ((~g28495));
assign g19196 = ((~II25423));
assign g21076 = ((~g20539));
assign g21881 = ((~g18492))|((~g19264))|((~g19278));
assign g30924 = (g30783&g22359);
assign g10558 = (g3366&g5150);
assign g8666 = (g7303&g7420);
assign g24451 = ((~g23644))|((~g3306));
assign gbuf50 = (g331);
assign g18837 = ((~g13998)&(~g12376));
assign g12970 = ((~g8523)&(~g8538)&(~g8551));
assign g22294 = ((~g20746));
assign g30651 = ((~g16265)&(~g30452));
assign g22558 = ((~II29116));
assign g30584 = ((~g30412)&(~g2611));
assign g8983 = ((~g6486));
assign g18838 = ((~g15248));
assign II18187 = ((~g7391));
assign g13714 = ((~g12453));
assign II29960 = ((~g22612));
assign II18130 = ((~g5547));
assign g4379 = ((~g1116));
assign g26854 = ((~II35011));
assign g12385 = ((~II19545));
assign g21006 = ((~g19828)&(~g17876));
assign II31706 = ((~g23836));
assign g6190 = ((~g2059));
assign g26538 = ((~g25458));
assign g20602 = ((~II27131));
assign II22989 = ((~g15296))|((~II22988));
assign g20673 = ((~II27264));
assign II14822 = ((~g1231));
assign gbuf118 = (g1309);
assign g25000 = (g24013)|(g24038);
assign g19014 = ((~II25105));
assign g22105 = ((~g21368)&(~g19664));
assign g13737 = ((~g13280));
assign g5714 = ((~g507));
assign II34662 = ((~g26174));
assign g23791 = ((~II31005));
assign II20802 = ((~g13160));
assign g26213 = (g25895&g9306);
assign II21554 = ((~g13074));
assign II36438 = ((~g27255));
assign g18923 = ((~g15582));
assign g5422 = ((~II13980));
assign g5991 = ((~g1651));
assign g22002 = ((~g21065))|((~g21711));
assign g25366 = ((~g24889));
assign g16252 = (g5813&g11899);
assign g13187 = ((~g9450));
assign g8102 = ((~g27));
assign II24207 = ((~g14102))|((~II24205));
assign g15467 = ((~II21726));
assign g18868 = ((~g14143)&(~g12419));
assign II29619 = ((~g21054));
assign g12306 = ((~g10598)&(~g10643)&(~g10674));
assign g29282 = ((~g28796));
assign g30733 = ((~II40487));
assign II35783 = ((~g26931));
assign II23904 = ((~g13561));
assign g27498 = ((~II35852));
assign g22353 = ((~II28913));
assign g27214 = ((~II35479));
assign g15033 = ((~g12030));
assign g21889 = ((~g19285)&(~g19316));
assign g16736 = ((~g14922)&(~g15065));
assign g26620 = ((~g25703));
assign g12518 = ((~g8655));
assign g29458 = ((~II38755));
assign g16513 = (g15065&g13724&g13764&g13797);
assign g8448 = (g6574&g1612);
assign g19178 = ((~g17718)&(~g15452));
assign g24833 = ((~g24245))|((~g24252));
assign g12915 = ((~g8955));
assign g15786 = ((~g12611))|((~g6369));
assign II25711 = ((~g2124))|((~II25710));
assign II24351 = ((~g14238))|((~g9356));
assign g28716 = (g28449&g19319);
assign II40191 = ((~g30360));
assign g27516 = (g23974&g27151);
assign g19070 = ((~g18583));
assign II13820 = ((~g797));
assign II30586 = ((~g23132));
assign g25249 = ((~g24821)&(~g23671));
assign II18055 = ((~g5668));
assign II22518 = ((~g13647));
assign II15354 = ((~g2574));
assign II16532 = ((~g7901));
assign g9883 = ((~II16880))|((~II16881));
assign II26505 = ((~g16693));
assign g13381 = ((~II20476));
assign II37474 = ((~g27762));
assign g13154 = ((~g9212));
assign g24951 = ((~II32709))|((~II32710));
assign II29632 = ((~g21061));
assign g17336 = ((~II23424));
assign II40444 = ((~g30591));
assign II31171 = ((~g23033));
assign II38518 = ((~g28783));
assign g25349 = ((~g24848));
assign g28695 = ((~II37632));
assign gbuf185 = (g2425);
assign II36882 = ((~g27987));
assign g22379 = ((~g20830));
assign g25856 = ((~II33700));
assign II40931 = ((~g30820));
assign II37757 = ((~g28512));
assign g24542 = (g19950&g18007&g23410);
assign g19924 = (g16551&g16924&g16529);
assign g24681 = ((~g24183)&(~g533));
assign g10123 = (g5473&g1116);
assign g22828 = ((~II29613));
assign II16338 = ((~g7015));
assign g26383 = (g4956&g25678);
assign g20011 = (g18063&g3113);
assign II41099 = ((~g30962));
assign g16725 = ((~II22741));
assign g18141 = ((~II24149))|((~II24150));
assign g27099 = (g22118&g26652);
assign g13989 = (g7661&g12894);
assign g24218 = ((~g16997)&(~g22264));
assign g28954 = ((~g26673)&(~g27241)&(~g28323));
assign II36909 = ((~g28006));
assign g16694 = ((~II22726));
assign g9121 = (g3774&g7760);
assign g7949 = ((~g165));
assign g24091 = ((~g22922))|((~g14438));
assign g27115 = (g5335&g26501);
assign g20322 = ((~g17327));
assign II33984 = ((~g25932));
assign g30801 = ((~g16237)&(~g30698));
assign g24920 = ((~II32660))|((~II32661));
assign g11662 = ((~g9534))|((~g3366));
assign g27124 = ((~g26410))|((~g5512));
assign II30738 = ((~g22067));
assign g27090 = (g23395&g26647);
assign gbuf74 = (g870);
assign g28500 = ((~g27794));
assign g25311 = ((~g24964)&(~g24029));
assign g22785 = ((~II29547));
assign g11351 = ((~II18305));
assign II30962 = ((~g22139));
assign g23330 = ((~g22186)&(~g22777));
assign II22676 = ((~g14630));
assign g18406 = ((~II24427))|((~II24428));
assign g30358 = ((~II39889));
assign g12463 = ((~g10730));
assign II24339 = ((~g6632))|((~II24338));
assign II40083 = ((~g30264));
assign II13131 = ((~g27));
assign g15847 = ((~g12611))|((~g6519));
assign g20556 = ((~II26993));
assign g26985 = (g14124&g26251);
assign II16296 = ((~g3306));
assign g28267 = ((~II37050));
assign g26944 = ((~g26374));
assign g20522 = ((~g16501))|((~g16515));
assign g12990 = (g8180&g10276);
assign g24219 = ((~g16998)&(~g22265));
assign g17942 = ((~II23982))|((~II23983));
assign II30233 = ((~g22833));
assign II32391 = ((~g17903))|((~g24034));
assign g30223 = (g30044&g9016);
assign g24456 = ((~g23803))|((~g3774));
assign gbuf157 = (g1946);
assign g10192 = (g3254&g4453);
assign II18332 = ((~g3566));
assign g19088 = (g18656&g14797&g16189&g13706);
assign g4433 = ((~g2255));
assign g15320 = (g7964&g12744);
assign g21488 = (g9857&g20451);
assign g26478 = (g5272&g25844);
assign g19032 = ((~II25159));
assign g24852 = ((~II32491))|((~II32492));
assign g5417 = ((~II13965));
assign g29137 = ((~II38154));
assign II25078 = ((~g15065));
assign II16056 = ((~g7606));
assign g13851 = (g7579&g12688);
assign g30087 = (g29840&g11120);
assign g18983 = ((~II25041));
assign II36314 = ((~g27575))|((~g15952));
assign g25814 = ((~II33652));
assign g22611 = ((~II29191));
assign g12476 = ((~g8622));
assign g8097 = ((~g2858));
assign g23022 = ((~g16968)&(~g21086));
assign g20998 = ((~II27549));
assign g18218 = ((~g14702))|((~g9928));
assign II25061 = ((~g14976));
assign g14767 = (g13245&g10765);
assign g28068 = ((~II36647));
assign g7779 = ((~g2395));
assign II33364 = ((~g25029));
assign II27200 = ((~g20479));
assign g21312 = (g9737&g20308);
assign g25363 = ((~g24862));
assign g24753 = ((~II32266))|((~II32267));
assign g21214 = ((~II27779));
assign g25463 = ((~II33289));
assign II33016 = ((~g25122));
assign II24253 = ((~g14520))|((~II24251));
assign g3365 = ((~g499));
assign II26282 = (g18188&g18089&g17991);
assign g19778 = (g18014&g16057);
assign II17429 = (g6901&g7338&g7146);
assign II15890 = ((~g3806));
assign II14571 = ((~g1145));
assign g4959 = ((~g1959));
assign g11559 = ((~II18653));
assign g19769 = (g17903&g16055);
assign II34916 = ((~g26240));
assign II27158 = ((~g20439));
assign g11213 = ((~II18139));
assign g26866 = (g5833&g26076);
assign g8996 = ((~II16312));
assign g17082 = (g7865&g15579);
assign g8549 = (g6519&g894);
assign II37197 = ((~g27903));
assign g22732 = (g18281&g21594);
assign g30933 = ((~g30755)&(~g30758));
assign II18866 = ((~g10875));
assign g26406 = (g5053&g25720);
assign g9793 = (g6980&g4049);
assign g23197 = ((~II30044));
assign II25897 = ((~g2147))|((~g18226));
assign g17582 = ((~II23670));
assign g26997 = (g22050&g26565);
assign g15920 = ((~g12657))|((~g6574));
assign g28298 = ((~II37143));
assign II37647 = ((~g28343));
assign g14614 = ((~g12293));
assign g7802 = ((~g2039));
assign g23115 = ((~g21708));
assign g11842 = ((~g11051));
assign II14009 = ((~g963));
assign g19111 = (g14936&g18772&g18796&g16433);
assign g28301 = ((~II37152));
assign g21453 = (g9941&g20434);
assign g7974 = ((~g3077));
assign II24613 = ((~g15978))|((~II24611));
assign g24093 = ((~g22922))|((~g14332));
assign II36915 = ((~g28007));
assign g13797 = ((~g12454));
assign g22970 = ((~II29736));
assign g17085 = ((~II23083))|((~II23084));
assign g30691 = ((~g13491)&(~g30355));
assign g13935 = ((~g11839));
assign g21647 = ((~II28174));
assign gbuf173 = (g2351);
assign g27715 = ((~II36156));
assign g23593 = (g22845&g20365);
assign g13687 = ((~g12460));
assign g23033 = ((~g21732))|((~g2746));
assign g12456 = ((~g8602));
assign g8430 = ((~g3198)&(~g8120)&(~g3194)&(~g3191));
assign g21007 = ((~g19829)&(~g15519));
assign g26970 = (g21976&g26544);
assign g30029 = ((~g29573)&(~g29962));
assign g22309 = (g1466&g21598);
assign g19345 = ((~II25732))|((~II25733));
assign g4740 = ((~g388));
assign g11899 = ((~g11148));
assign g5856 = ((~II14306));
assign g12312 = ((~II19479));
assign II17081 = ((~g3338));
assign g8575 = ((~II15779));
assign g19329 = ((~II25711))|((~II25712));
assign II38245 = ((~g28920));
assign g24546 = ((~g23898)&(~g22770));
assign II16225 = ((~g6042));
assign g27007 = (g23360&g26580);
assign g17616 = (g6626&g16041);
assign g8478 = ((~II15680));
assign g19555 = (g8001&g17243);
assign II25308 = ((~g16867));
assign gbuf119 = (g1312);
assign g20620 = ((~II27185));
assign g10839 = ((~g5798)&(~g5846)&(~g5882));
assign II25762 = ((~g79))|((~II25761));
assign g18115 = ((~II24132))|((~II24133));
assign II20441 = ((~g9027));
assign g15852 = (g7878&g11642);
assign g25808 = ((~II33646));
assign g10924 = ((~II17807));
assign g20278 = ((~g17237));
assign g8443 = ((~II15645));
assign g18152 = (g5218&g15701);
assign g25282 = (g24648&g8748);
assign g17058 = ((~II23046))|((~II23047));
assign g26308 = ((~II34266));
assign g30480 = ((~II40054));
assign g11702 = ((~g9676))|((~g3522));
assign g21046 = ((~g19887)&(~g15650));
assign g5621 = ((~g3161));
assign g30876 = ((~II40880));
assign II37203 = ((~g27912));
assign II23999 = ((~g15074));
assign g29402 = ((~g29077));
assign g15785 = ((~g12565))|((~g6314));
assign II13098 = ((~g2637));
assign II40587 = ((~g30629))|((~g30622));
assign g27269 = ((~g26997)&(~g26293));
assign g20911 = ((~g19667)&(~g17528));
assign g26761 = (g26154&g22257);
assign II35841 = ((~g26807));
assign g23684 = ((~II30844));
assign g29291 = ((~g28817));
assign g29528 = (g28750&g29369);
assign g30342 = ((~II39853));
assign II15616 = ((~g6838));
assign g13443 = ((~II20628));
assign gbuf33 = (g284);
assign II14378 = ((~g3234));
assign g21164 = ((~II27727));
assign g13061 = ((~g9676))|((~g6980));
assign g20136 = (g17878&g9423);
assign g21175 = (g20178&g12366);
assign g24862 = ((~II32527))|((~II32528));
assign g19661 = (g653&g18823);
assign g12099 = ((~g10305)&(~g10382)&(~g10446));
assign II24601 = ((~g6890))|((~g14135));
assign g18270 = ((~II24264))|((~II24265));
assign g24596 = (g771&g23887);
assign II13149 = ((~g45));
assign II25344 = ((~g17847));
assign II29513 = ((~g21019));
assign gbuf198 = (g2619);
assign g27839 = ((~II36307));
assign g27850 = ((~g27501)&(~g14650));
assign II40985 = ((~g30792));
assign II23639 = ((~g15900));
assign g29918 = ((~g29744)&(~g22367));
assign II24481 = ((~g15993));
assign g27018 = (g22005&g26586);
assign g11721 = ((~g9534))|((~g3366));
assign g25209 = ((~g24749)&(~g23554));
assign g16995 = ((~II22946))|((~II22947));
assign g4058 = ((~g1534));
assign g21501 = (g20522)|(g16867)|(g14071);
assign II30254 = ((~g22659));
assign g24777 = (g12876&g24130);
assign g15830 = ((~g13310))|((~g12392));
assign II16101 = ((~g3878));
assign gbuf17 = (g2851);
assign g23089 = (g21806)|(g21799);
assign II32509 = ((~g17815))|((~g24070));
assign g8784 = (g7391&g8242);
assign II24150 = ((~g14408))|((~II24148));
assign g12833 = ((~II19894));
assign II17486 = ((~g3900));
assign g23429 = ((~g23107));
assign g10725 = ((~g3710))|((~g7230));
assign II22759 = ((~g14703));
assign II30639 = ((~g22038));
assign g15396 = ((~II21658));
assign g5849 = ((~II14295));
assign g13118 = ((~g9822))|((~g7230));
assign g11776 = ((~g10943));
assign g30364 = (g30211&g8452);
assign g29538 = (g29210&g29376);
assign g29072 = ((~g9342))|((~g28595));
assign g12759 = ((~II19823));
assign II40973 = ((~g30784));
assign II30791 = ((~g22846))|((~II30790));
assign g27046 = (g22093&g26612);
assign II37994 = ((~g28556));
assign II29209 = ((~g20911));
assign II40886 = ((~g30819));
assign II23266 = ((~g14413))|((~II23264));
assign g24691 = (g24103)|(g20866);
assign g8275 = ((~II15493));
assign g16458 = (g5996&g12173);
assign g29924 = ((~g29710)&(~g22367));
assign II24745 = ((~g14486))|((~II24743));
assign g10583 = (g3650&g1982);
assign II18686 = ((~g9932));
assign g9133 = (g3462&g7796);
assign II30194 = ((~g22685));
assign g16282 = (g5835&g11918);
assign g25342 = (g5851&g24600);
assign g26800 = ((~g26163)&(~g25457));
assign g4515 = ((~g1119));
assign II24317 = ((~g6832))|((~g14217));
assign g19602 = (g633&g18785);
assign g17114 = (g8242&g15638);
assign g29522 = (g27735&g29363);
assign g25599 = ((~II33424));
assign g8249 = ((~II15429));
assign g11890 = ((~g9890)&(~g10010)&(~g10103));
assign II28065 = ((~g19957));
assign II15794 = ((~g3338));
assign g20610 = ((~II27155));
assign II18076 = ((~g3566));
assign g9774 = (g6678&g4023);
assign g23587 = ((~II30673));
assign g12481 = ((~g8627));
assign g29206 = ((~g28909)&(~g28459));
assign g16017 = (g12130&g10862);
assign g17301 = (g8097&g15994);
assign g26202 = ((~II34118));
assign II25320 = ((~g16924));
assign g11287 = ((~II18235));
assign g24315 = ((~II31619));
assign g27154 = ((~II35347));
assign g12440 = ((~II19598));
assign g4970 = ((~g2097));
assign g20658 = ((~g20198))|((~g3410));
assign g12412 = ((~II19560));
assign g7826 = ((~g2987));
assign II40664 = ((~g30636));
assign g28640 = ((~g27928));
assign II34012 = ((~g25938));
assign II28148 = ((~g19987));
assign g12146 = ((~g10369)&(~g10436)&(~g10496));
assign g29581 = ((~g29406)&(~g17065));
assign g5390 = ((~II13896));
assign II36441 = ((~g27256));
assign g10183 = (g7426&g4444);
assign g16131 = ((~g12871));
assign g20567 = ((~II27026));
assign II40435 = ((~g30585));
assign g29266 = ((~g28741));
assign g11370 = ((~II18326));
assign g19125 = ((~II25320));
assign g18928 = ((~g15606));
assign II17737 = ((~g6000));
assign g27360 = ((~II35678));
assign g22987 = ((~g21646)&(~g21068));
assign II33909 = ((~g25886));
assign g23602 = ((~II30704));
assign g8613 = (g6945&g7349);
assign II39539 = ((~g29911))|((~g29913));
assign g17993 = ((~g14016));
assign g17710 = ((~II23794));
assign g19678 = (g4185&g17479);
assign II25495 = (g17158)|(g17137)|(g17115);
assign g12101 = ((~g11444));
assign g13550 = ((~g12657))|((~g3566));
assign II13904 = ((~g358));
assign g27052 = (g4885&g26358);
assign g25950 = ((~g24574)&(~g24580));
assign g20063 = (g5382&g18569);
assign g11692 = ((~g9676))|((~g3522));
assign g30930 = ((~g30735)&(~g30744));
assign g22715 = ((~II29399));
assign II24368 = ((~g15990));
assign II21577 = ((~g12981));
assign g25143 = ((~II32907));
assign II36781 = ((~g15151))|((~II36779));
assign g23715 = (g17937&g23006);
assign g21731 = (g3710&g20535);
assign g18089 = ((~g14355));
assign g12245 = ((~g10495)&(~g10557)&(~g10604));
assign g5084 = ((~g1962));
assign g23205 = ((~II30068));
assign g30804 = ((~II40664));
assign g4480 = ((~g707));
assign g9676 = (g7788&g6145&g1224);
assign g18708 = ((~g14863));
assign g26003 = ((~II33861));
assign II14882 = ((~g1786));
assign g17758 = ((~II23833));
assign II19862 = ((~g10725));
assign g23768 = (g4570&g22629);
assign g19816 = (g2026&g18900);
assign g16289 = (g5853&g11929);
assign g16138 = (g5641&g11820);
assign g7999 = ((~g485));
assign g9893 = (g6448&g420);
assign g16134 = (g5363&g11818);
assign II28876 = ((~g21238));
assign g4685 = ((~g1724));
assign II17849 = ((~g8103));
assign g22945 = ((~II29724));
assign g13525 = ((~g12657))|((~g3566));
assign g22033 = ((~g21301)&(~g19560));
assign g28555 = ((~II37488));
assign g30783 = ((~g30618)&(~g22387));
assign g28336 = (g27896&g20810);
assign g11995 = ((~g11303));
assign g10498 = (g3462&g5041);
assign g25990 = ((~II33822));
assign II18683 = ((~g9733));
assign g28705 = ((~II37662));
assign g26683 = ((~II34656));
assign g29502 = (g29350&g8912);
assign g8176 = ((~g2845));
assign II24280 = ((~g13918))|((~II24278));
assign II14544 = ((~g1041));
assign g15897 = ((~g12657))|((~g6783));
assign II17846 = ((~g8107));
assign II38028 = ((~g28584));
assign g29654 = ((~II39080));
assign II22884 = ((~g13370))|((~g15661));
assign g23679 = (g4304&g22567);
assign II38632 = ((~g29298));
assign g29818 = (g29732&g22293);
assign g24463 = ((~g23923))|((~g3338));
assign II25004 = ((~g14459));
assign g11386 = ((~II18344));
assign g7724 = ((~g2389));
assign II33831 = ((~g25982));
assign II30272 = ((~g22797));
assign g23264 = ((~II30245));
assign g10451 = (g3618&g4945);
assign II32443 = ((~g18014))|((~g24054));
assign g11629 = ((~II18813));
assign II33737 = ((~g24476));
assign g12292 = ((~g10584)&(~g10625)&(~g10660));
assign g15664 = ((~g12565))|((~g6314));
assign II33882 = ((~g25364));
assign g29388 = ((~g29023));
assign g7329 = ((~g2734));
assign II29249 = ((~g20923));
assign g11965 = ((~g10094)&(~g10184)&(~g10272));
assign II34118 = ((~g25605));
assign g8755 = (g3494&g8004);
assign g29724 = ((~g29500));
assign g12223 = ((~g8427));
assign g28350 = ((~g15604)&(~g28057));
assign g26364 = ((~II34327));
assign g28746 = ((~g15046)&(~g28441));
assign g8570 = (g3566&g1591);
assign II24452 = ((~g6142))|((~g14450));
assign g11873 = ((~g9794)&(~g9921)&(~g10058));
assign g22165 = ((~g21444)&(~g19773));
assign g10522 = (g3678&g5089);
assign II33561 = ((~g25047));
assign g18224 = ((~g14592));
assign g23845 = ((~II31085));
assign II36948 = ((~g27976));
assign II27110 = ((~g19622));
assign g13740 = (g6636&g12547);
assign g25157 = ((~II32949));
assign II27243 = ((~g19335));
assign g15480 = ((~II21739));
assign g30658 = ((~g16312)&(~g30462));
assign II34026 = ((~g25892));
assign II14049 = ((~g870));
assign g28080 = (g27604&g10130);
assign II35777 = ((~g27119));
assign II21256 = ((~g11647));
assign II28210 = ((~g20537));
assign II25682 = ((~g70))|((~II25681));
assign g28701 = ((~II37650));
assign II30519 = ((~g22942));
assign g28273 = ((~II37068));
assign g10012 = (g3306&g423);
assign II27182 = ((~g20458));
assign g8395 = (g6519&g912);
assign g27323 = ((~g27071)&(~g26423));
assign g8719 = ((~II15925));
assign g5975 = ((~g2333));
assign g5397 = ((~II13907));
assign g26961 = (g13907&g26175);
assign II39347 = ((~g29732))|((~g29728));
assign g29120 = ((~II38128));
assign II29484 = ((~g21903));
assign g3960 = ((~g861));
assign g28897 = (g14016&g28641);
assign g19571 = (g8153&g17294);
assign g16749 = ((~g15782));
assign g24106 = ((~g22428));
assign g28485 = (g18453&g28178);
assign g25978 = (g24836&g13850);
assign g21775 = ((~g20198))|((~g6369));
assign g26592 = ((~g13851)&(~g25300));
assign g17165 = ((~II23208))|((~II23209));
assign g8161 = ((~g2218));
assign g20357 = ((~g16743)&(~g16974));
assign g16050 = (g5590&g11764);
assign II38606 = ((~g29039));
assign g13952 = (g7643&g12881);
assign II17936 = ((~g6314));
assign II18969 = ((~g8726));
assign II18163 = ((~g6574));
assign g20946 = ((~g19733)&(~g17654));
assign g20937 = ((~g19717)&(~g17620));
assign II18737 = ((~g8910));
assign g25745 = ((~g20866)&(~g24440));
assign g17949 = (g4970&g15569);
assign II21822 = ((~g13106));
assign g12353 = (g7852&g8915);
assign g28081 = ((~II36684));
assign g7785 = ((~g1010));
assign g18755 = ((~g13871)&(~g12274));
assign g29415 = ((~II38626));
assign g27235 = ((~II35542));
assign g21035 = ((~g19874)&(~g18013));
assign g18120 = ((~g14115));
assign g9090 = (g7391&g2641);
assign II17925 = ((~g7976));
assign II13849 = ((~g1486));
assign g22939 = ((~g21877))|((~g21875))|((~g21873));
assign g7685 = ((~g1091));
assign g12054 = ((~g11386));
assign II34433 = ((~g25271));
assign g5912 = ((~g2160));
assign g12952 = ((~g10252)&(~g6626));
assign g7389 = ((~g2185));
assign g18876 = ((~g15418));
assign g30836 = ((~II40760));
assign II24387 = ((~g6421))|((~g13974));
assign g23377 = ((~g21968))|((~g22308));
assign g28036 = (g14541&g27535);
assign II36942 = ((~g27905));
assign II14496 = ((~g3226));
assign g6713 = ((~II14819));
assign g9302 = (g6232&g7993);
assign g25140 = ((~II32898));
assign II31868 = ((~g23719));
assign g29696 = ((~II39142));
assign g15851 = ((~g12711))|((~g7085));
assign g19665 = (g4133&g17457);
assign II21340 = ((~g11779));
assign gbuf65 = (g543);
assign II40787 = ((~g30809));
assign g13332 = ((~g11481)&(~g8045)&(~g11190)&(~g7880));
assign g30775 = ((~II40588))|((~II40589));
assign g3338 = ((~II13169));
assign g28305 = ((~II37164));
assign II36404 = ((~g27450));
assign g27571 = ((~g26869))|((~g56));
assign II19195 = ((~g8726));
assign g18552 = ((~g16154));
assign g23161 = ((~II29936));
assign g22272 = (g21742&g12282);
assign II37961 = ((~g28501));
assign g8350 = (g6574&g1594);
assign g5605 = ((~g3182));
assign g16104 = (g12235&g10946);
assign g8659 = ((~II15853));
assign II31931 = ((~g23725));
assign g20389 = ((~g17531));
assign g24176 = ((~g22600));
assign II15429 = ((~g2833));
assign II40167 = ((~g30456));
assign g18912 = ((~g15537));
assign II23163 = ((~g13857))|((~II23161));
assign g10457 = (g7053&g4959);
assign II22718 = ((~g14657));
assign II40441 = ((~g30586));
assign g21605 = (g19067)|(g19524)|(g16529);
assign II31853 = ((~g23676));
assign II34755 = ((~g26206));
assign g30120 = ((~II39625));
assign g29133 = ((~II38142));
assign g24328 = ((~II31658));
assign g11928 = ((~g10008)&(~g10102)&(~g10192));
assign II30868 = ((~g22881))|((~g14194));
assign g22949 = ((~g21665));
assign g23112 = ((~g21700));
assign g29008 = ((~g9174))|((~g28540));
assign g3995 = ((~g3064));
assign g27467 = ((~II35809));
assign g15691 = ((~II21942));
assign g20904 = ((~g19896));
assign g29784 = ((~g29484)&(~g29236));
assign g12213 = ((~g10453)&(~g10516)&(~g10572));
assign g30109 = (g29857&g11411);
assign g19146 = (g17191&g16788);
assign g7560 = ((~g2526));
assign g21244 = (g19578)|(g16697)|(g14776);
assign g25274 = ((~g24912));
assign g13495 = ((~g12611))|((~g3410));
assign g4289 = ((~g2082));
assign II37775 = ((~g28540));
assign g12524 = ((~g10315)&(~g10393)&(~g10455));
assign g16908 = (g7838&g15032);
assign gbuf26 = (g276);
assign g29660 = ((~g29578));
assign g10251 = (g7230&g4555);
assign g21339 = (g9326&g20336);
assign g19730 = (g653&g17573);
assign g18958 = ((~g15714));
assign II28365 = (g20280)|(g18652)|(g18649);
assign g23214 = ((~II30095));
assign g13139 = ((~g9968))|((~g7488));
assign g10519 = (g7053&g5084);
assign II29194 = ((~g20902));
assign g8421 = ((~II15623));
assign II33529 = ((~g25041));
assign II36156 = ((~g27586));
assign g21157 = (g5809&g19291);
assign II23504 = ((~g15848));
assign g18950 = ((~g15688));
assign g12994 = ((~g8542)&(~g8555)&(~g8564));
assign g29313 = ((~g28717)&(~g19117));
assign g24441 = (g14737&g15981&g24168);
assign g12782 = ((~g8836));
assign g29952 = (g29784&g28959);
assign II18004 = ((~g3410));
assign II26497 = (g18212)|(g18115)|(g18030);
assign g28734 = ((~g28525));
assign g4304 = ((~g2247));
assign g18469 = ((~g14497));
assign II36693 = ((~g27320));
assign g24623 = ((~g24183)&(~g529));
assign II27149 = ((~g19893));
assign g13175 = ((~g8725)&(~g8762)&(~g8783));
assign g15133 = ((~II21446));
assign g19749 = ((~II26182));
assign II36933 = ((~g28049));
assign g16183 = (g12235&g11014);
assign II24363 = ((~g14525))|((~II24361));
assign II20820 = ((~g13171));
assign g29571 = ((~g28710)&(~g29176));
assign g27295 = ((~g27029)&(~g26362));
assign g25401 = ((~g24823));
assign II25099 = ((~g19000));
assign II15912 = ((~g3878));
assign II40997 = ((~g30797));
assign II18572 = ((~g8931));
assign g30982 = ((~II41120));
assign g17215 = ((~g15904)&(~g14642));
assign g14291 = ((~g12050));
assign g23272 = ((~II30269));
assign g5890 = ((~g88));
assign g13011 = ((~II20062));
assign g27028 = (g22050&g26599);
assign g8636 = (g7391&g7535);
assign g30649 = ((~g16253)&(~g30449));
assign g18880 = ((~g15443));
assign g18652 = (g14797&g13657&g13677&g16243);
assign II25243 = ((~g17227));
assign g30407 = (g30134&g10991);
assign g23485 = ((~II30531));
assign g10642 = (g3834&g5280);
assign g29550 = (g29222&g29385);
assign II30032 = ((~g22672));
assign g30283 = ((~g16431)&(~g30118));
assign g10003 = ((~II16966))|((~II16967));
assign II39909 = ((~g30291));
assign g30187 = ((~g30023));
assign II21626 = ((~g11693));
assign g22555 = (g13895&g21415);
assign II16684 = ((~g6486));
assign II32178 = ((~g24237));
assign II34779 = ((~g26308));
assign g26693 = ((~II34686));
assign g19654 = (g4098&g17433);
assign g20718 = ((~g20228))|((~g3566));
assign g5224 = ((~g2794));
assign g6170 = ((~g3098));
assign II26695 = (g18670&g18692&g16142);
assign II37796 = ((~g28634));
assign II21165 = ((~g13110));
assign g11802 = ((~g10991));
assign g8859 = ((~II16107));
assign g11883 = ((~g11120));
assign g6116 = ((~II14631));
assign II40032 = ((~g30254));
assign g24286 = ((~II31532));
assign g10101 = (g3254&g4329);
assign g11385 = ((~II18341));
assign II25666 = ((~g18474))|((~II25664));
assign II39469 = ((~g29935));
assign g28970 = (g14322&g28651);
assign g27314 = ((~g27056)&(~g26404));
assign g23105 = ((~II29852));
assign g29148 = ((~II38187));
assign g19846 = (g1358&g18914);
assign g24612 = ((~II32198));
assign g11347 = (g6232&g213);
assign g25265 = ((~g24878)&(~g23852));
assign g15048 = ((~g12045));
assign g12004 = ((~g11324));
assign g24253 = (g21995&g11370);
assign g10850 = ((~II17701));
assign g23970 = ((~g22887))|((~g14119));
assign g18648 = (g14811&g14976&g16201&g13791);
assign II37394 = ((~g27718));
assign II25351 = ((~g17959));
assign II25126 = ((~g16858));
assign g4263 = ((~g1411));
assign II23860 = ((~g15932));
assign II40524 = ((~g30690));
assign II38386 = ((~g28734));
assign g17715 = (g4581&g15379);
assign g26840 = ((~II34983));
assign g26553 = ((~g13816)&(~g25282));
assign g20227 = (g13714&g13756&II26661);
assign II36283 = ((~g27408));
assign II14027 = ((~g182));
assign g4912 = ((~II13680));
assign g24898 = (g24060&g18931);
assign II22786 = ((~g14725));
assign g28065 = (g27608&g10070);
assign g8022 = ((~g2930));
assign g27927 = ((~II36390));
assign g24144 = ((~g22506));
assign g24365 = ((~II31769));
assign g24842 = ((~II32461))|((~II32462));
assign II36711 = ((~g27325));
assign g18206 = ((~II24206))|((~II24207));
assign g7540 = ((~g1506));
assign g30442 = (g30155&g11111);
assign g17797 = (g4731&g15449);
assign g26374 = ((~g25964)&(~g24503));
assign II30215 = ((~g22766));
assign g19726 = (g16847&g6131);
assign g30132 = (g30068&g20776);
assign g26619 = ((~g25700));
assign g26209 = ((~g25296));
assign II24464 = ((~g14360))|((~g9453));
assign g4538 = ((~g1546));
assign g24559 = (g79&g23448);
assign g4809 = ((~g1690));
assign g4979 = ((~g2115));
assign g4788 = ((~g1396));
assign g5263 = ((~g2466));
assign g17221 = ((~g4848)&(~g14618));
assign g18435 = ((~g14359));
assign II16630 = ((~g6057));
assign g3460 = ((~II13182));
assign g5241 = ((~g1297));
assign g11278 = ((~II18226));
assign g5825 = ((~g1684));
assign II40122 = ((~g30443));
assign g28098 = (g27604&g10214);
assign g24388 = ((~II31838));
assign g24605 = ((~II32189));
assign g12289 = ((~g8469));
assign g24497 = ((~g23734)&(~g22638));
assign II27399 = ((~g19390));
assign g28137 = ((~g27566));
assign g25216 = ((~g24757)&(~g23565));
assign g13423 = ((~II20568));
assign II17363 = ((~g3806));
assign g26731 = ((~II34800));
assign g29253 = ((~II38360));
assign g29305 = ((~II38450));
assign g12252 = ((~g8443));
assign g4592 = ((~g361));
assign II16117 = ((~g5473));
assign g22041 = ((~g21308)&(~g19568));
assign g26877 = ((~g26140)&(~g22319));
assign g19451 = ((~II25881))|((~II25882));
assign II38421 = ((~g28740));
assign g16370 = (g5917&g12003);
assign g9115 = (g3618&g7742);
assign II31493 = ((~g23587));
assign II37629 = ((~g28369));
assign g28171 = (g27349&g10898);
assign g23871 = ((~II31127));
assign g19007 = (g14976&g13687&g13714&g13756);
assign g16488 = ((~II22566));
assign g24552 = (g18598&g23107&g23410);
assign g10056 = (g7162&g4257);
assign g28979 = ((~II37946));
assign g4250 = ((~g1107));
assign g14130 = (g7724&g12960);
assign g29082 = ((~II38049));
assign II38683 = ((~g29308));
assign II35545 = ((~g26964));
assign g22503 = ((~II29049));
assign g20429 = ((~g17679));
assign g15638 = ((~g12373));
assign g29260 = (g28863&g8934);
assign g20269 = ((~g17230));
assign g27527 = ((~g26759)&(~g19087));
assign II29500 = ((~g21015));
assign g27021 = (g23335&g26589);
assign II23695 = ((~g15870));
assign g9782 = (II16826&II16827);
assign g8336 = ((~II15538));
assign g15672 = ((~II21923));
assign g23284 = ((~II30305));
assign II16166 = ((~g6713));
assign II19996 = (g9795&g9711&g9595&g9471);
assign II40805 = ((~g30767));
assign II26664 = ((~g17847));
assign g9407 = ((~g5945));
assign g9519 = (g6314&g8194);
assign g26576 = ((~II34535));
assign II32982 = ((~g24612));
assign g22744 = ((~II29468));
assign II29168 = ((~g20775));
assign II16247 = ((~g5422));
assign g26260 = (g25254&g17649);
assign g20732 = ((~II27321));
assign g17173 = ((~II23226))|((~II23227));
assign g28990 = ((~g28667)&(~g16457));
assign II33520 = ((~g25062));
assign g23413 = ((~g17694)&(~g22654));
assign II13110 = ((~g8));
assign g23826 = ((~II31050));
assign g18679 = ((~g14811));
assign II26231 = ((~g18401));
assign g17439 = ((~II23527));
assign g25949 = ((~g24565)&(~g24573));
assign g11265 = ((~II18211));
assign g18441 = ((~II24465))|((~II24466));
assign g29992 = (g12441&g29909);
assign g20766 = ((~II27355));
assign g26178 = ((~II34080));
assign g23238 = ((~II30167));
assign g24747 = (g9427&g24099);
assign II24966 = ((~g14863));
assign g22851 = ((~g16113)&(~g20850)&(~g21278));
assign g21390 = (g9174&g20385);
assign II15623 = ((~g7085));
assign II32156 = ((~g24225));
assign g13389 = ((~II20486));
assign II18370 = ((~g4093))|((~II18368));
assign II30041 = ((~g22706));
assign II38148 = ((~g29074));
assign g28224 = ((~II36921));
assign II32409 = ((~g18131))|((~g24037));
assign II38710 = ((~g29408));
assign g23945 = ((~g4456)&(~g13565)&(~g23009));
assign g21113 = ((~II27672));
assign g13163 = ((~g9273));
assign g22336 = ((~g20216)&(~g21818));
assign II37260 = ((~g28179));
assign II40925 = ((~g30752));
assign II40307 = ((~g30500));
assign g29709 = ((~g29583)&(~g1909));
assign g23567 = (g8233&g22440);
assign II20794 = ((~g13111));
assign g5107 = ((~g2448));
assign g12369 = ((~g10680)&(~g10707)&(~g10724));
assign g7334 = ((~II14957));
assign II25325 = ((~g16954));
assign g28652 = ((~g27994));
assign g26832 = ((~II34967));
assign g10980 = ((~II17881));
assign g24478 = (g23545&g21119&g21227);
assign g20088 = (g16836&g3147);
assign g4447 = ((~g2801));
assign II36407 = ((~g27581));
assign II13221 = ((~g2241));
assign g4038 = ((~g859));
assign g6019 = ((~g1471));
assign gbuf200 = (g2587);
assign II25198 = ((~g16878));
assign g10169 = (g7085&g4424);
assign g20942 = ((~II27488));
assign g19222 = (g18195)|(g18441);
assign g23135 = ((~g21229)&(~g19449));
assign II16759 = ((~g3462));
assign II31799 = ((~g23532));
assign g4766 = ((~g736));
assign II35319 = ((~g26183));
assign g14459 = ((~g12151));
assign II32548 = ((~g23906))|((~II32546));
assign g9725 = (g6783&g3975);
assign II13275 = ((~g2848));
assign g28966 = (g28625&g9481);
assign II37901 = ((~g28529));
assign g8852 = ((~II16098));
assign g21489 = (g15366&g20452);
assign g3978 = ((~g1554));
assign g18744 = ((~g14936));
assign g13190 = ((~g9481));
assign II33879 = ((~g25488));
assign II39124 = ((~g29606));
assign g22200 = ((~g21553)&(~g19883));
assign g30322 = ((~II39809));
assign g5917 = ((~g2315));
assign g30022 = ((~g29547)&(~g29955));
assign II32922 = ((~g24577));
assign g9127 = (g3306&g7782);
assign g13053 = ((~g9968))|((~g7488));
assign g11830 = ((~g9647)&(~g9773)&(~g9901));
assign g4339 = ((~II13433));
assign II39376 = ((~g29768))|((~II39375));
assign II33870 = ((~g25797));
assign g30812 = ((~II40688));
assign g17856 = ((~II23917));
assign g15631 = ((~II21884));
assign g30488 = ((~II40066));
assign g26702 = ((~II34713));
assign g27779 = (g5760&g27367);
assign g11727 = ((~g9822))|((~g3678));
assign g30055 = ((~g29965)&(~g13326));
assign II27137 = ((~g19596));
assign g5952 = ((~II14416));
assign g19647 = (g2020&g18813);
assign g26712 = ((~II34743));
assign g15017 = ((~g12009));
assign g10886 = ((~g5889));
assign II32081 = ((~g24178));
assign g22262 = ((~g20690));
assign g10932 = ((~II17819));
assign II39385 = ((~g29718))|((~II39384));
assign II38122 = ((~g28421));
assign gbuf150 = (g1931);
assign II13990 = ((~g2463));
assign g19753 = (g2033&g18860);
assign II36582 = ((~g27291));
assign g20542 = ((~g16523))|((~g16546));
assign g22300 = ((~II28876));
assign g20470 = ((~II26913));
assign g10397 = (g7358&g4836);
assign II13215 = ((~g2009));
assign II32561 = ((~g24081))|((~II32559));
assign g17734 = (g4611&g15393);
assign g10219 = (g6980&g4523);
assign g27751 = ((~g25400))|((~g27455));
assign g24902 = (g18469&g23874);
assign g28844 = (g27850&g28582);
assign g5306 = ((~g2102));
assign g5416 = ((~II13962));
assign g21064 = ((~II27621));
assign g17342 = ((~II23430));
assign II40490 = ((~g30679));
assign g8514 = ((~g6139));
assign g24513 = ((~g15425)&(~g23843));
assign g8265 = ((~II15463));
assign g24561 = (g18598&g23429&g19975);
assign g28778 = ((~g28464)&(~g27963));
assign II35297 = ((~g26199));
assign g24392 = ((~II31850));
assign g28412 = (g7812&g27879);
assign g27454 = ((~g26783)&(~g25196));
assign II36423 = ((~g27466));
assign II37356 = ((~g27824))|((~g27811));
assign II34680 = ((~g26294));
assign g19681 = ((~g16974));
assign II18317 = ((~g3410));
assign g21227 = ((~g18414)&(~g18485)&(~g20295));
assign II37608 = ((~g28455));
assign g22266 = ((~g20694));
assign g13537 = ((~g12565))|((~g3254));
assign II22875 = ((~g14966));
assign g27427 = (g2072&g27139);
assign g25082 = ((~g23428)&(~g22207));
assign II18335 = ((~g6783));
assign g13435 = ((~II20604));
assign II34353 = ((~g25927));
assign II20601 = ((~g13321));
assign g25128 = (g17051&g24115&g13614);
assign II19482 = ((~g10500));
assign g12843 = ((~g8879));
assign II33807 = ((~g25588));
assign II36585 = ((~g27292));
assign II38007 = ((~g28556));
assign g17048 = (g7845&g15493);
assign gbuf190 = (g2447);
assign II18506 = ((~g8699));
assign II18417 = ((~g6574));
assign g23473 = ((~II30519));
assign g10096 = ((~II17066));
assign g10676 = ((~g3398))|((~g6678));
assign g27748 = ((~g27632));
assign g29624 = (g29254&g11407);
assign gbuf114 = (g1229);
assign g27705 = ((~II36126));
assign II14900 = ((~g2211));
assign II31298 = ((~g22280));
assign g26679 = ((~II34644));
assign g27562 = ((~II35968));
assign g5677 = (g331&g366);
assign II20649 = ((~g13344));
assign II16018 = ((~g6058));
assign II14113 = ((~g1012));
assign II25429 = ((~g18975));
assign g8284 = ((~II15499));
assign g13905 = (g7925&g12847);
assign g16033 = (g5546&g11748);
assign g15274 = ((~g11875));
assign g16836 = ((~g15818));
assign g12808 = ((~II19869));
assign g22360 = ((~g20822));
assign g14390 = ((~g12971));
assign g15323 = ((~g12242));
assign g28480 = (g18297&g27977);
assign g5378 = ((~g2933));
assign g5182 = ((~g1965));
assign g5731 = ((~g1192));
assign g11813 = ((~g11004));
assign II32335 = ((~g23997))|((~II32333));
assign g22310 = ((~g20776));
assign g18519 = ((~g13741));
assign g10087 = ((~II17051));
assign g21099 = ((~II27658));
assign II22813 = ((~g13601));
assign g10021 = ((~II16993));
assign g28164 = ((~g27440));
assign g9065 = (g3494&g1176);
assign II31244 = ((~g22687));
assign g22998 = ((~g21458));
assign g28041 = ((~g27376));
assign II30134 = ((~g22559));
assign g13404 = ((~g8183)&(~g11332)&(~g7928)&(~g7880));
assign g19628 = (g653&g18807);
assign g20981 = ((~g19795)&(~g17795));
assign II40462 = ((~g30670));
assign II21415 = ((~g11854));
assign g29823 = ((~g29663));
assign g13093 = ((~g9822))|((~g7230));
assign g24909 = (g23726)|(g23142);
assign II15800 = ((~g3494));
assign g24993 = ((~g23521));
assign g21566 = ((~II28100));
assign g26345 = (g25261&g17850);
assign II22640 = ((~g14650));
assign II39770 = ((~g30063));
assign g19943 = (g7562&g18976);
assign II13943 = ((~g2418));
assign g27181 = (g16570&g26508&g13614);
assign II14624 = ((~g1155));
assign g25942 = ((~g24805));
assign II32913 = ((~g24586));
assign II21720 = ((~g11701));
assign II24475 = ((~g6184))|((~II24474));
assign g29117 = ((~II38119));
assign II34689 = ((~g26433));
assign g24525 = ((~g15495)&(~g23866));
assign II13320 = ((~g2864));
assign g18843 = ((~g15271));
assign g17724 = ((~g13886));
assign g9613 = ((~g5876));
assign II13119 = ((~g17));
assign g6832 = ((~g2033));
assign II32526 = ((~g18038))|((~g24078));
assign g13397 = ((~II20500));
assign g28393 = ((~II37330));
assign g26738 = ((~II34821));
assign g19552 = (g16829&g6048);
assign g22691 = ((~II29345));
assign II39466 = ((~g29934));
assign g19718 = (g4295&g17545);
assign g6031 = ((~II14502));
assign g28406 = ((~g27824)&(~g22344));
assign g19848 = (g1365&g18916);
assign g21102 = ((~g19081));
assign g5772 = ((~g1193));
assign g29958 = (g29783&g29027);
assign g28055 = ((~II36618));
assign II34071 = ((~g25212));
assign g7519 = ((~II15019));
assign g27567 = ((~g4809)&(~g26891));
assign g18352 = ((~g16082)&(~g14249));
assign g22288 = ((~g20144)&(~g21805));
assign II29030 = ((~g20683));
assign g19318 = ((~II25682))|((~II25683));
assign II40275 = ((~g30375));
assign g25228 = ((~g24776)&(~g23590));
assign g26587 = ((~g25599));
assign g11904 = ((~g11157));
assign II16200 = ((~g7303));
assign II28184 = ((~g19103));
assign g17465 = ((~II23553));
assign g29357 = ((~g29129)&(~g17100));
assign g25119 = ((~II32847));
assign g24533 = ((~g23864)&(~g22738));
assign g5818 = ((~g1194));
assign II15526 = ((~g6314));
assign g15577 = (g5113&g13241);
assign g30713 = ((~II40429));
assign g27475 = ((~II35817));
assign II40257 = ((~g30488));
assign g4671 = ((~g1563));
assign g5286 = ((~g2797));
assign g28377 = ((~II37284));
assign II18392 = ((~g6369));
assign g19605 = (g3951&g17357);
assign g27485 = ((~g26928)&(~g24638));
assign g29249 = ((~II38352));
assign g10401 = (g3722&g4851);
assign II27041 = ((~g19237));
assign g10225 = (g5512&g4541);
assign g17464 = (g4153&g15139);
assign g20576 = ((~II27053));
assign g28117 = ((~II36776));
assign g10540 = (g7488&g5135);
assign g13071 = ((~g9534))|((~g6678));
assign II38199 = ((~g29100));
assign g26041 = ((~g25475)&(~g24855));
assign g15144 = ((~g12109));
assign g19152 = ((~g5378))|((~g18884));
assign g20487 = ((~g18308))|((~g2026));
assign g19058 = ((~II25237));
assign g30334 = (g30203&g8347);
assign g16070 = (g12187&g10921);
assign g26819 = ((~II34946));
assign g7009 = ((~g1352));
assign g30704 = ((~g14040)&(~g30392));
assign II26416 = (g18553&g18491&g18431);
assign II37252 = ((~g28200));
assign g11028 = ((~II17939));
assign g17670 = ((~II23754));
assign g3878 = ((~II13242));
assign II35849 = ((~g26776));
assign II33545 = ((~g25045));
assign g5719 = ((~g909));
assign g24281 = ((~II31517));
assign g23394 = ((~g18572))|((~g22887));
assign g23292 = ((~II30329));
assign g15403 = (g4623&g12786);
assign g21142 = (g20000&g20020);
assign II18016 = ((~g5720));
assign g8329 = (g6232&g231);
assign g28367 = ((~g15769)&(~g28122));
assign g8708 = ((~II15912));
assign II24677 = ((~g6305))|((~g14637));
assign g10080 = (g7085&g4307);
assign II13999 = ((~g276));
assign II39791 = ((~g30126));
assign g27737 = (g27558&g16832);
assign g27150 = ((~II35341));
assign II31130 = ((~g22184));
assign g28877 = ((~II37846));
assign g25231 = ((~g24780)&(~g23599));
assign g13233 = ((~g9898));
assign g29397 = ((~g29065));
assign g29327 = ((~II38502));
assign g5954 = ((~g192));
assign II27733 = (g19277&g19451&g19416);
assign II18250 = ((~g3566));
assign g11496 = ((~II18464));
assign g19761 = (g2766&g18865);
assign g8934 = ((~II16228));
assign II37614 = ((~g28580));
assign g13340 = (g5727&g11294);
assign g29242 = (g9737&g28826);
assign g13942 = ((~g11843));
assign II18692 = ((~g10935));
assign g21181 = (g20242&g12373);
assign g9911 = (g5473&g1104);
assign g14486 = ((~g12171));
assign g10210 = (g5473&g4512);
assign g22281 = (g21782&g12296);
assign g13339 = ((~II20410));
assign g7581 = ((~g1496));
assign g26558 = ((~g25515));
assign g19952 = (g2760&g18987);
assign g8866 = ((~II16120));
assign g29332 = (g29080&g29019);
assign g23553 = ((~II30607));
assign II25174 = ((~g18971));
assign g19907 = (g17954&g18390&II26357);
assign II16697 = ((~g6713));
assign g30096 = (g29844&g11268);
assign g27083 = (g22093&g26640);
assign g29577 = ((~g28714)&(~g29186));
assign g5145 = ((~g584));
assign g5811 = ((~g801));
assign II17027 = ((~g3650));
assign g10865 = ((~g6131));
assign g28294 = ((~II37131));
assign g8560 = ((~g3554))|((~g3522));
assign II26528 = (g18656&g14837&g13657);
assign g16841 = ((~g15021)&(~g12607));
assign g22582 = ((~II29142));
assign g6145 = ((~II14660));
assign g27061 = (g23372&g26627);
assign II14897 = ((~g2211));
assign g21554 = ((~II28084));
assign g18699 = ((~g14849));
assign g11809 = ((~g10999));
assign g10078 = (g6838&g4301);
assign g30849 = ((~II40799));
assign g21793 = ((~g19515)&(~g18237)&(~g14431));
assign II20500 = ((~g11007));
assign g8014 = ((~II15308));
assign g28348 = ((~g15594)&(~g28050));
assign g23155 = ((~II29918));
assign g12321 = ((~II19488));
assign g8254 = ((~g3063));
assign g4861 = ((~II13655));
assign g16445 = (g5808&g13381);
assign g22517 = (g21895&g12608);
assign II33469 = ((~g24498));
assign g5163 = ((~g1300));
assign g26765 = (g26399&g19265);
assign g28826 = ((~II37787));
assign g23999 = ((~g22922))|((~g14234));
assign g23776 = (g18074&g23021);
assign g18453 = ((~g14472));
assign II23715 = ((~g15931));
assign g30743 = (g30610&g22283);
assign g20247 = (g14936&g18772&g16325&g16371);
assign II17203 = ((~g6115));
assign g8267 = ((~II15469));
assign II21813 = ((~g13104));
assign g5934 = ((~g942));
assign g10325 = (g3722&g4711);
assign g29932 = ((~II39398));
assign g18337 = ((~g15757));
assign g21863 = ((~g18212))|((~g19205))|((~g19213));
assign g19748 = (g4398&g17610);
assign g12083 = ((~g10293)&(~g10371)&(~g10438));
assign g11734 = ((~g10843));
assign g27733 = (g27513&g16785);
assign g19559 = (g8059&g17255);
assign g26639 = ((~g25784));
assign g21452 = (g6427&g19749);
assign g11741 = ((~g10880));
assign g19211 = (g18441)|(g18497);
assign II40116 = ((~g30408));
assign II38752 = ((~g29276));
assign g14115 = ((~II21083));
assign g21720 = ((~g14256))|((~g15177))|((~g19871))|((~g19842));
assign g30537 = ((~II40191));
assign g23265 = ((~II30248));
assign g6025 = ((~g2264));
assign g18997 = (g13541&g16278);
assign g30479 = ((~II40051));
assign g20416 = ((~g17627));
assign g8832 = ((~II16062));
assign g15175 = ((~g12139));
assign II39325 = ((~g29713))|((~II39323));
assign gbuf161 = (g1908);
assign g28145 = ((~g27629)&(~g17001));
assign g8150 = ((~g1525));
assign g29370 = ((~g28928));
assign g18346 = ((~II24352))|((~II24353));
assign g29687 = ((~g29572)&(~g29344));
assign g4174 = ((~g1789));
assign II25117 = ((~g18988));
assign g22701 = (g18174&g21561);
assign g8552 = (g6783&g1579);
assign II24522 = ((~g14234))|((~II24520));
assign g26079 = ((~g25445))|((~g25413))|((~g25301));
assign g28936 = (g28619&g9384);
assign g10433 = (g3338&g602);
assign II37787 = ((~g28595));
assign g27900 = ((~g6087)&(~g27632)&(~g25338));
assign g13913 = (g7623&g12850);
assign II15553 = ((~g3566));
assign g10818 = ((~g5740)&(~g5787)&(~g5826));
assign g16018 = (g6149&g11741);
assign g29552 = ((~g29130)&(~g29411));
assign g12561 = ((~II19733));
assign g26465 = ((~II34425));
assign g26087 = ((~g6068)&(~g24183)&(~g25319));
assign g25031 = ((~g23694))|((~g5473));
assign g30341 = ((~g14328)&(~g30226));
assign g19181 = (g17729)|(g17979);
assign II22671 = ((~g14691));
assign g19637 = (g4055&g17410);
assign g10392 = (g7015&g1822);
assign g16298 = (g520&g11936);
assign II36462 = ((~g27259));
assign g29815 = (g29727&g20662);
assign II38740 = ((~g29288));
assign II33006 = ((~g24957));
assign g26594 = ((~g25620));
assign II18476 = ((~g8791));
assign g13625 = (g6173&g12476);
assign g20094 = (g13677&g13706&II26528);
assign II13169 = ((~g550));
assign g26423 = (g5107&g25749);
assign II32479 = ((~g17927))|((~II32478));
assign g19731 = (g646&g18853);
assign II18429 = ((~g7085));
assign II32410 = ((~g18131))|((~II32409));
assign g17100 = (g3722&g10754&g14493);
assign g16386 = (g5933&g12037);
assign g20599 = ((~II27122));
assign g28467 = ((~II37426));
assign g17779 = ((~II23854));
assign g7697 = ((~g2388));
assign g10075 = (g7358&g4292);
assign II25691 = ((~g753))|((~II25690));
assign g14724 = (g7861&g13117);
assign g10015 = ((~g5292));
assign g26743 = ((~II34836));
assign g30495 = (g30179&g11422);
assign II27897 = ((~g19149));
assign g10628 = (g7358&g5260);
assign II30191 = ((~g22715));
assign g4298 = ((~g2231));
assign g23335 = ((~g23096))|((~g23083));
assign g8635 = (g3650&g7354);
assign g25749 = ((~II33580));
assign II29238 = ((~g20919));
assign g28228 = ((~II36933));
assign g23582 = (g3975&g22464);
assign g21736 = ((~g20164))|((~g6232));
assign g8828 = ((~II16056));
assign II19865 = ((~g10354));
assign g30858 = ((~II40826));
assign g24584 = ((~II32146));
assign g12789 = ((~g8340)&(~g8395)&(~g8437));
assign II32708 = ((~g23892))|((~g14402));
assign g17451 = ((~II23539));
assign g5121 = ((~g2664));
assign g21779 = ((~g20545)&(~g18567));
assign II18139 = ((~g6643));
assign g9427 = ((~g5645));
assign g27167 = ((~g26474));
assign g24027 = ((~g22922))|((~g14139));
assign II31490 = ((~g23569));
assign g27679 = (g26782&g11386);
assign g14630 = ((~II21241));
assign g19195 = (g17942)|(g18212);
assign g10682 = (g3774&g5335);
assign II30269 = ((~g22769));
assign g6425 = ((~g974));
assign g8180 = ((~g3071));
assign g25717 = ((~II33545));
assign g25132 = ((~II32874));
assign g30579 = ((~II40291));
assign II39933 = ((~g30298));
assign g23716 = (g22886&g20432);
assign g21353 = (g9326&g20351);
assign g14006 = (g7670&g12914);
assign II24372 = ((~g14454))|((~g9310));
assign g10645 = (g3834&g5289);
assign II25159 = ((~g18913));
assign II13680 = ((~g813));
assign g21447 = (g15274&g20430);
assign g28855 = ((~g28409));
assign g8272 = ((~II15484));
assign g16632 = ((~g15981)&(~g15971)&(~g14711));
assign g17523 = ((~II23611));
assign II23235 = ((~g14291))|((~II23233));
assign g21010 = ((~g19840)&(~g17901));
assign g14525 = ((~g12195));
assign g15160 = (g4313&g13174);
assign g26796 = ((~II34921));
assign g12104 = ((~g11453));
assign g21049 = (g20016&g14079&g14165);
assign II28488 = ((~g21495));
assign g30268 = ((~g16382)&(~g30102));
assign II19576 = ((~g10683));
assign g7909 = ((~II15226));
assign g5592 = ((~g515));
assign g26080 = (g25950&g21164);
assign g28178 = ((~g27518));
assign g5832 = ((~g1921));
assign g15442 = (g2714&g12804);
assign g30668 = ((~g16381)&(~g30478));
assign II29013 = ((~g21764));
assign g21580 = ((~g20067));
assign g19479 = ((~g16733));
assign g30901 = ((~II40955));
assign II14917 = ((~g1312));
assign II36513 = ((~g27272));
assign g24323 = ((~II31643));
assign g23042 = ((~g21778)&(~g21143));
assign g24125 = ((~g22467));
assign g29923 = ((~II39360))|((~II39361));
assign II21852 = ((~g11716));
assign g17046 = ((~II23019))|((~II23020));
assign II39982 = ((~g30305));
assign II30689 = ((~g22054));
assign II16538 = ((~g3306));
assign g24407 = ((~II31895));
assign II23460 = ((~g13501));
assign II21772 = ((~g13097));
assign II28582 = (g19141&g21133&g21116);
assign g22396 = ((~g21219))|((~g14529))|((~g10714));
assign g23742 = (g23119)|(g21920);
assign g16089 = (g984&g11787);
assign g14558 = ((~g12217));
assign g28425 = ((~g16133)&(~g28188));
assign gbuf95 = (g1074);
assign g28215 = ((~II36894));
assign g27838 = ((~II36301))|((~II36302));
assign g27188 = ((~g26091)&(~g25388));
assign g16953 = (g7482&g15144);
assign g30908 = ((~II40976));
assign II24291 = ((~g13895))|((~II24290));
assign g15034 = ((~II21389));
assign II40572 = ((~g30588))|((~II40571));
assign g13104 = ((~g9676))|((~g7162));
assign g4746 = ((~g580));
assign g13089 = ((~g9534))|((~g6912));
assign g20562 = ((~II27011));
assign II15276 = ((~g2935))|((~g2938));
assign g27372 = (g2133&g27064);
assign gbuf136 = (g1731);
assign g28358 = ((~g15700)&(~g28094));
assign II21420 = ((~g13166));
assign g29691 = ((~II39127));
assign g24261 = ((~II31457));
assign g27990 = ((~g27367));
assign g29795 = ((~II39237));
assign g5735 = ((~g1476));
assign g19530 = ((~g16817));
assign g19061 = ((~II25246));
assign II28755 = ((~g13541))|((~II28753));
assign g28285 = ((~II37104));
assign g30083 = (g29835&g11048);
assign g11120 = ((~II18034));
assign g30452 = (g30163&g11166);
assign g10710 = (g3806&g2694);
assign II30941 = ((~g22131));
assign g15475 = (g4928&g13220);
assign g27012 = ((~g26668)&(~g21931));
assign g29171 = ((~II38250));
assign g12446 = ((~g8605)&(~g10773));
assign g11766 = ((~g10886));
assign II34815 = ((~g26250));
assign II24752 = ((~g7455))|((~II24751));
assign g12908 = (g7899&g10004);
assign II32696 = ((~g23858))|((~II32695));
assign g22804 = (g2920&g21655);
assign g18988 = ((~II25054));
assign II34761 = ((~g26245));
assign g15814 = ((~II22063))|((~II22064));
assign II17928 = ((~g8031));
assign g27147 = ((~g23458)&(~g26054));
assign g22381 = ((~g21211))|((~g14442))|((~g10694));
assign gbuf128 = (g1835);
assign g25354 = ((~II33188));
assign II39895 = ((~g30287));
assign g28900 = ((~II37871));
assign g29081 = ((~II38046));
assign g19001 = ((~g14071));
assign g8873 = ((~g4955));
assign g28312 = ((~II37185));
assign II19872 = ((~g8317));
assign g6188 = ((~g1904));
assign g23249 = ((~II30200));
assign g7961 = ((~II15267));
assign g13298 = ((~g10235));
assign g10290 = (g6678&g4617);
assign II17786 = ((~g7193));
assign g14001 = ((~g12849));
assign II24632 = ((~g7009))|((~g14467));
assign g30052 = ((~II39550));
assign g15246 = (g4475&g13186);
assign g28727 = ((~g28489));
assign g7353 = ((~g1140));
assign g8794 = ((~II15998));
assign g13042 = (g8100&g10601);
assign II21787 = ((~g11707));
assign II14499 = ((~g3214));
assign II34728 = ((~g26264));
assign II15345 = ((~g1862));
assign g27449 = ((~g26837));
assign g5398 = ((~II13910));
assign g24989 = (g23983)|(g24004);
assign g29915 = ((~II39340))|((~II39341));
assign g5427 = ((~II13993));
assign II34710 = ((~g26214));
assign g6058 = ((~II14553));
assign g11867 = ((~g11095));
assign II32940 = ((~g24562));
assign II18220 = ((~g6232));
assign g21636 = ((~g20473)&(~g6513));
assign II18689 = ((~g10231));
assign g4476 = ((~g576));
assign g9105 = (g3462&g7712);
assign g14212 = (g7736&g12972);
assign II37575 = ((~g28527));
assign g9957 = (g6838&g4197);
assign g30674 = ((~g16414)&(~g30492));
assign II15308 = ((~g1880));
assign g13705 = (g12776&g8673);
assign g29390 = ((~g29032));
assign II22881 = ((~g13622));
assign g29369 = ((~g28925));
assign II32609 = ((~g24090))|((~II32607));
assign g30014 = ((~g29526)&(~g29947));
assign g22328 = ((~II28896));
assign II33652 = ((~g25072));
assign g7346 = ((~g97));
assign g19015 = ((~II25108));
assign g27586 = ((~II36008));
assign g13069 = ((~g9968))|((~g7426));
assign g25015 = ((~g23694))|((~g6713));
assign II35491 = ((~g26956));
assign g14342 = ((~g12967));
assign II38220 = ((~g29102));
assign g23849 = (g22771&g17868);
assign g20368 = ((~g17457));
assign II35686 = ((~g27131));
assign g10424 = ((~g7910));
assign g27855 = ((~g6087)&(~g27632)&(~g25385));
assign g10207 = (g6519&g4501);
assign II16176 = ((~g7936));
assign g11055 = ((~II17972));
assign II40478 = ((~g30675));
assign g16290 = (g5854&g11930);
assign g4516 = ((~g1125));
assign II31778 = ((~g23794));
assign g30374 = (g30211&g8475);
assign g8745 = ((~II15935));
assign g21094 = ((~g19952)&(~g18404));
assign II19932 = ((~g10763));
assign g12551 = ((~g8700));
assign g18902 = ((~g15502));
assign g16571 = (g15913)|(g14691);
assign g29216 = ((~g28940)&(~g28472));
assign II35803 = ((~g26803));
assign g24304 = ((~II31586));
assign g5027 = ((~g581));
assign g28364 = ((~g15740)&(~g28112));
assign g30729 = ((~II40475));
assign g12222 = ((~g8424));
assign g28280 = ((~II37089));
assign II40185 = ((~g30346));
assign g25240 = ((~g24798)&(~g23622));
assign g19128 = ((~g16708))|((~g16728));
assign g5808 = ((~g509));
assign g24881 = (g24047&g18912);
assign II16559 = ((~g5512));
assign g23624 = (g17741&g22989);
assign II16169 = ((~g5405));
assign g30387 = (g30229&g8888);
assign II35530 = ((~g26910));
assign II22663 = ((~g14711));
assign II31757 = ((~g23744));
assign g8810 = ((~II16018));
assign II40850 = ((~g30724));
assign g30179 = ((~g30021));
assign g7927 = ((~g3076));
assign g16011 = ((~g12651));
assign II34428 = ((~g25931));
assign g13347 = ((~g10409));
assign g6573 = ((~II14783));
assign II30988 = ((~g22145));
assign g26578 = ((~g25573));
assign g12020 = ((~g11341));
assign g8521 = (g3410&g951);
assign g27328 = ((~g27080)&(~g26437));
assign g19097 = (g13657&g16243&II25280);
assign g16536 = ((~g15873))|((~g2896));
assign II17206 = ((~g3650));
assign g19785 = (g2026&g18878);
assign g25647 = ((~II33472));
assign g8809 = ((~II16015));
assign g12494 = (g7833&g9134);
assign g13264 = ((~g10096));
assign g28455 = ((~II37410));
assign g20992 = ((~g19805)&(~g15470));
assign g26327 = ((~g25958)&(~g24493));
assign II19591 = ((~g8900));
assign II36093 = ((~g27514));
assign g5800 = ((~II14246));
assign g27342 = ((~g27098)&(~g26473));
assign g20950 = ((~g19742)&(~g17674));
assign II36786 = ((~g27343));
assign II30508 = ((~g23047));
assign g16042 = ((~g12765));
assign g11781 = ((~g9442)&(~g9522)&(~g9633));
assign g28355 = ((~g15671)&(~g28080));
assign II21548 = ((~g11684));
assign II27209 = ((~g20485));
assign g13172 = ((~g9335));
assign g21427 = ((~II27972));
assign II31417 = ((~g22578));
assign g9390 = ((~II16593));
assign g29970 = (g29764&g12178);
assign II32994 = ((~g24865));
assign g13893 = ((~g8580))|((~g12463));
assign II32997 = ((~g24903));
assign II29093 = ((~g21791));
assign II38038 = ((~g28346));
assign II16714 = ((~g5512));
assign II35673 = ((~g27123));
assign II40152 = ((~g30359));
assign g30720 = ((~II40450));
assign II17753 = ((~g6943));
assign II36752 = ((~g27335));
assign II24582 = ((~g15996));
assign g18629 = (g13764&g13819&II24738);
assign g25762 = ((~II33593));
assign g14228 = (g7745&g12979);
assign g16835 = ((~g15717)&(~g12966));
assign g24357 = ((~II31745));
assign g8305 = ((~g3805));
assign g5683 = ((~g789));
assign II37149 = ((~g28093));
assign II22998 = ((~g9187))|((~g13872));
assign g26968 = (g6305&g26542);
assign g15339 = (g4655&g13200);
assign g4348 = ((~g704));
assign II14644 = ((~g3142));
assign II21381 = ((~g13157));
assign g6041 = ((~II14516));
assign II32092 = ((~g23418));
assign g16417 = (g5759&g13356);
assign II18320 = ((~g6519));
assign g5323 = ((~g2798));
assign II38437 = ((~g28736));
assign g26244 = (g25903&g9387);
assign g21029 = ((~g19864)&(~g15592));
assign II21479 = ((~g13035));
assign g10855 = ((~g5847)&(~g5883)&(~g5919));
assign II34180 = ((~g25240));
assign g29129 = ((~g28385)&(~g27790));
assign II20414 = ((~g8575));
assign II27194 = ((~g20484));
assign g27799 = ((~II36250));
assign II14928 = ((~g1931));
assign g26346 = (g25911&g9727);
assign g24033 = ((~II31253));
assign g26980 = (g23360&g26554);
assign g10441 = (g3494&g4919);
assign II15593 = ((~g6519));
assign g24893 = ((~g23486));
assign g6637 = ((~g5));
assign g16528 = ((~II22611));
assign gbuf180 = (g2359);
assign g28730 = ((~g28470));
assign g20450 = ((~g17776));
assign g4070 = ((~g1557));
assign g24234 = ((~g22289)&(~g21157));
assign II29326 = ((~g20952));
assign g19249 = ((~II25510));
assign II28323 = (g20227)|(g20211)|(g20183);
assign g29473 = (g21508&g29269);
assign g10822 = ((~g5748)&(~g5797)&(~g5845));
assign g12478 = ((~g10749));
assign g23893 = (g22966&g9933);
assign g8535 = (g6519&g885);
assign g20978 = ((~g19785)&(~g17774));
assign g20697 = ((~II27288));
assign g21646 = ((~g20058)&(~g14194)&(~g14280));
assign II14945 = ((~g2480));
assign II15511 = ((~g8014));
assign II38674 = ((~g29177));
assign g12271 = ((~g10538)&(~g10597)&(~g10642));
assign g10367 = (g3366&g4754);
assign g24756 = ((~g16089)&(~g24211));
assign g4090 = ((~II13320));
assign g24700 = (g17217&g24168);
assign II20390 = ((~g10821));
assign g24950 = ((~g23710));
assign g15823 = ((~g12611))|((~g6519));
assign g9886 = ((~g7149));
assign g6051 = ((~II14532));
assign II35136 = ((~g26660));
assign g13157 = ((~g9229));
assign g8827 = ((~II16053));
assign g24489 = ((~g23674)&(~g22596));
assign g14098 = (g7709&g12944);
assign II15185 = ((~g2978))|((~II15183));
assign II37017 = ((~g28113));
assign g19987 = ((~II26437));
assign g13229 = ((~II20278));
assign g22641 = ((~II29249));
assign II17834 = ((~g7976));
assign g28739 = ((~g28429)&(~g27915));
assign g26445 = (g5176&g25787);
assign g26393 = ((~II34353));
assign g11603 = ((~II18777));
assign g26770 = (g26059&g19287);
assign g20682 = ((~g19160)&(~g10024));
assign g7349 = ((~g1167));
assign g23059 = ((~g14490)&(~g14412)&(~g21162));
assign g25046 = ((~g23748))|((~g5512));
assign g17634 = (g4447&g15317);
assign g9075 = (g6448&g7643);
assign II14868 = ((~g1237));
assign gbuf176 = (g2527);
assign II33304 = ((~g25004));
assign g21678 = ((~II28206));
assign II25801 = ((~g83))|((~II25800));
assign g10170 = (g6838&g4427);
assign g17542 = (g4286&g15225);
assign II33961 = ((~g25357));
assign II24445 = ((~g9507))|((~II24443));
assign g26777 = (g26066&g19305);
assign g26215 = ((~II34143));
assign g27121 = ((~g26367))|((~g5473));
assign II28009 = ((~g20473));
assign g23178 = ((~II29987));
assign g16243 = ((~g13033));
assign g28944 = (g28625&g9404);
assign II40643 = ((~g30568));
assign g21000 = ((~g19817)&(~g17854));
assign g14520 = ((~g12184));
assign g8980 = ((~II16296));
assign g23835 = ((~II31065));
assign g25041 = ((~g23923))|((~g6643));
assign g4383 = ((~g1392));
assign II20619 = ((~g13366));
assign g27696 = ((~II36099));
assign II16110 = ((~g5404));
assign g27265 = ((~g26993)&(~g26288));
assign II19886 = ((~g10706));
assign II35933 = ((~g26950));
assign g20648 = ((~g20164))|((~g3254));
assign g19250 = (g17729)|(g17807);
assign g10280 = (g6448&g4595);
assign g29110 = ((~g28656)&(~g17031));
assign II24594 = ((~g6438))|((~g14139));
assign g18430 = ((~g16020)&(~g14352));
assign g19806 = (g4629&g17738);
assign g15655 = ((~II21908));
assign g18961 = ((~g15726));
assign g10910 = ((~II17789));
assign g16934 = ((~II22881));
assign II18827 = ((~g10936));
assign g7776 = ((~g1009));
assign II36749 = ((~g27334));
assign g19255 = (g14366)|(g16523);
assign g19820 = (g18131&g16093);
assign g28886 = ((~g28659)&(~g16277));
assign g27559 = ((~II35961));
assign g21974 = ((~g20938)&(~g10340));
assign II29921 = ((~g23078));
assign g29155 = ((~II38208));
assign g16423 = (g5772&g13361);
assign II18638 = ((~g8826));
assign g20439 = ((~II26868));
assign II30023 = ((~g22550));
assign g20057 = (g18290)|(g18195)|(II26491);
assign g13857 = ((~g11760));
assign g16965 = ((~II22901))|((~II22902));
assign II38822 = ((~g15933))|((~II38820));
assign II40772 = ((~g30804));
assign II40988 = ((~g30793));
assign g30013 = ((~g29525)&(~g29946));
assign II19733 = ((~g8726));
assign g28299 = ((~II37146));
assign g25393 = ((~g24866));
assign gbuf79 = (g1141);
assign II15326 = ((~g3117));
assign g12460 = ((~II19642));
assign g30127 = (g30065&g20719);
assign g23165 = ((~II29948));
assign g25937 = ((~g24763));
assign g11428 = ((~II18392));
assign g16420 = (g5961&g12086);
assign g22621 = ((~II29209));
assign g21843 = ((~g13619)&(~g19155));
assign II18854 = ((~g10854));
assign II19533 = ((~g10631));
assign g30352 = (g30211&g8414);
assign g12198 = ((~II19374));
assign II25848 = ((~g18358))|((~II25846));
assign g12269 = ((~g10533)&(~g10592)&(~g10637));
assign g17345 = ((~II23433));
assign II18845 = ((~g10911));
assign g28251 = ((~II37002));
assign II37297 = ((~g27814))|((~II37295));
assign g5221 = ((~g2792));
assign II23338 = ((~g15721));
assign g4614 = ((~g715));
assign g14099 = ((~II21075));
assign II34321 = ((~g25928));
assign II27155 = ((~g20395));
assign II36224 = ((~g27589));
assign gbuf145 = (g1776);
assign g20093 = (g13657&g13677&g13750&II26525);
assign g24245 = (g19417)|(g22402);
assign II29369 = ((~g20967));
assign II26171 = ((~g17594));
assign g19335 = ((~II25728));
assign II19569 = ((~g10653));
assign g20690 = ((~II27281));
assign g26601 = ((~g25643));
assign g18727 = ((~g14966));
assign g10906 = ((~g5924));
assign g21254 = (g20318&g14910);
assign II38282 = ((~g28941));
assign gbuf51 = (g545);
assign II25477 = (g17024)|(g17000)|(g16992);
assign g30215 = ((~II39674));
assign II40420 = ((~g30578));
assign g21807 = (g16527)|(g19063)|(g19007)|(II28330);
assign g19541 = (g16913&g16764&g14811);
assign g28064 = ((~II36639));
assign II40568 = ((~g30701));
assign g19051 = ((~II25216));
assign g27865 = ((~g6087)&(~g27632)&(~g25370));
assign g24577 = ((~II32129));
assign g10362 = (g3338&g4743);
assign g29138 = ((~II38157));
assign II27176 = ((~g20469));
assign g20885 = ((~g19865));
assign II23559 = ((~g15869));
assign II34165 = ((~g25236));
assign g11719 = ((~g9822))|((~g3678));
assign g9749 = ((~II16793));
assign g26472 = ((~g16615))|((~g25195));
assign g24529 = (g19933&g17896&g23403);
assign II40811 = ((~g30772));
assign g16867 = ((~g13589));
assign II18817 = ((~g9067));
assign g30635 = ((~g16108)&(~g30407));
assign II25213 = ((~g18993));
assign g4555 = ((~g2088));
assign g25235 = ((~g24790)&(~g23606));
assign g20025 = ((~II26469));
assign g22108 = ((~g21789))|((~g21801));
assign II33507 = ((~g25058));
assign II30014 = ((~g22786));
assign g28015 = (g14472&g27518);
assign II32251 = ((~g23919));
assign II29525 = ((~g21023));
assign g16154 = ((~g12194));
assign g19951 = ((~II26407));
assign II18716 = ((~g8944));
assign II25228 = ((~g18937));
assign gbuf8 = (g2824);
assign g13398 = ((~g10542));
assign g28324 = (g27810&g20659);
assign II36612 = ((~g27298));
assign II29395 = ((~g20976));
assign II27278 = ((~g19369));
assign gbuf207 = (g2642);
assign II40634 = ((~g30571));
assign II32725 = ((~g23913))|((~II32724));
assign g5970 = ((~g1648));
assign g24772 = (g15618&g24124);
assign g18313 = ((~II24318))|((~II24319));
assign g28106 = ((~II36749));
assign g25988 = ((~II33816));
assign II24188 = ((~g13958))|((~II24186));
assign g9773 = (g6912&g4020);
assign II36099 = ((~g27515));
assign g15198 = ((~II21488));
assign g20282 = (g14849&g18728&g13687&g16302);
assign g29518 = (g28728&g29360);
assign g12898 = ((~g9407)&(~g9342));
assign g18169 = (g7527&g15714);
assign g5900 = ((~g933));
assign II26913 = ((~g17270));
assign g28156 = ((~g27410));
assign g22216 = ((~g21635)&(~g19944));
assign g19107 = (g17223&g16616);
assign g21402 = (g9427&g20398);
assign gbuf27 = (g405);
assign II13959 = ((~g1754));
assign II24417 = ((~g15366))|((~II24415));
assign g20876 = ((~g19585)&(~g17353));
assign g18854 = ((~g15329));
assign g18998 = ((~II25078));
assign g13201 = ((~g9607));
assign II27920 = ((~g19154));
assign g10379 = (g6945&g1276);
assign g13220 = ((~g9787));
assign g30541 = ((~II40203));
assign g30082 = (g29829&g11036);
assign g6945 = ((~II14868));
assign g29765 = ((~g13492)&(~g29465));
assign g25409 = ((~g24808));
assign g30752 = ((~II40534));
assign II30857 = ((~g22105));
assign II25645 = ((~g18190))|((~II25643));
assign g29489 = (g21580&g29296);
assign II23219 = ((~g13903))|((~II23217));
assign g19827 = (g2720&g18904);
assign g29468 = (g29343&g19490);
assign gbuf20 = (g3129);
assign II34734 = ((~g26407));
assign II13801 = ((~g2195));
assign II19833 = ((~g8726));
assign g30642 = ((~g16199)&(~g30440));
assign g22599 = ((~II29177));
assign g18947 = ((~g15675));
assign g13409 = ((~II20526));
assign g5355 = ((~g1425));
assign g22153 = ((~g21423)&(~g19755));
assign g20153 = ((~g16536)&(~g7583));
assign gbuf42 = (g367);
assign II33382 = ((~g25016));
assign g27484 = ((~g26855));
assign g27035 = (g23377&g26606);
assign g13252 = ((~II20305));
assign g5150 = ((~g722));
assign g22830 = (g14541&g21671);
assign g11502 = ((~II18482));
assign g15794 = ((~II22044));
assign II21806 = ((~g13103));
assign g5008 = ((~g2661));
assign g16858 = ((~II22836));
assign g27843 = ((~II36311));
assign g12090 = ((~g10297)&(~g10373)&(~g10439));
assign II16258 = ((~g3306));
assign g19944 = (g3028&g18258);
assign g13234 = ((~II20283));
assign II19829 = ((~g10631));
assign g18603 = ((~II24695))|((~II24696));
assign g22682 = (g2040&g21550);
assign g29744 = ((~g29583)&(~g24641));
assign II23982 = ((~g14292))|((~II23981));
assign g10596 = (g3834&g5218);
assign g21865 = ((~g18424))|((~g19210))|((~g19221));
assign g9150 = ((~g5893));
assign II26639 = (g18656&g18670&g16142);
assign II19777 = ((~g10735));
assign II15866 = ((~g3878));
assign g29057 = ((~II38014));
assign II29496 = ((~g21011));
assign g24480 = ((~g23617)&(~g23659));
assign g17824 = (g4766&g15471);
assign II36897 = ((~g28005));
assign g19091 = ((~II25272));
assign g30594 = ((~g6119)&(~g30412)&(~g25419));
assign g23850 = (g23139)|(g20647);
assign g11315 = ((~II18265));
assign g26886 = ((~II35083));
assign g28374 = ((~II37277));
assign II17768 = ((~g8031));
assign g5005 = ((~g2650));
assign g29168 = ((~II38245));
assign g15856 = ((~g12565))|((~g6232));
assign g27784 = ((~II36221));
assign II25050 = ((~g14601));
assign II31598 = ((~g23574));
assign g12452 = ((~II19628));
assign II24648 = ((~g9795))|((~II24646));
assign g30481 = (g30179&g11351);
assign g19566 = (g8129&g17278);
assign g29616 = ((~g13969)&(~g29259));
assign g22104 = ((~g21367)&(~g19663));
assign g22083 = ((~g21774))|((~g21787));
assign g21156 = (g19290&g19276&II27717);
assign g4437 = ((~g2492));
assign g16431 = (g5975&g12117);
assign g4688 = ((~g1750));
assign II34207 = ((~g25969));
assign g21271 = ((~II27822));
assign g20005 = ((~g18124));
assign g25071 = ((~g23984))|((~g7053));
assign g22048 = ((~g21314)&(~g19575));
assign g27349 = ((~g27126));
assign g17874 = (g4870&g15510);
assign g11647 = ((~g9079)&(~g9094)&(~g9103));
assign II23926 = ((~g15074));
assign g26352 = (g25919&g9749);
assign g24781 = (g12916&g24133);
assign g8029 = ((~g3083));
assign g6632 = ((~g2720));
assign g20002 = ((~II26444));
assign g19030 = ((~II25153));
assign g18096 = ((~II24111))|((~II24112));
assign g27922 = (g4112&g27416);
assign g13391 = ((~II20490));
assign g13261 = ((~g10070));
assign g30436 = (g30134&g11079);
assign II40432 = ((~g30582));
assign II30278 = ((~g22691));
assign g16647 = ((~II22690));
assign g13214 = ((~g9752));
assign g11822 = ((~g9632)&(~g9760)&(~g9888));
assign II39945 = ((~g30302));
assign g19457 = ((~II25904));
assign g29032 = ((~II37991));
assign g22673 = ((~II29313));
assign g29186 = (g29063&g20769);
assign g9453 = ((~g5717));
assign g7638 = ((~g2546));
assign g29968 = (g29765&g12119);
assign II35975 = ((~g27094))|((~II35974));
assign II24567 = ((~g9595))|((~II24565));
assign g29276 = ((~II38401));
assign II17975 = ((~g7265));
assign II38866 = ((~g29179));
assign g10568 = (g6945&g1294);
assign g25095 = ((~g23786));
assign g20965 = ((~g19761)&(~g17717));
assign g21399 = ((~II27942));
assign g6630 = ((~g1668));
assign II25867 = ((~g18573))|((~II25865));
assign g29861 = ((~g29677));
assign g25305 = ((~g24880));
assign g20164 = ((~II26612));
assign g20819 = ((~II27408));
assign g5403 = ((~II13925));
assign g21302 = (g9374&g20290);
assign g29075 = ((~II38038));
assign II29019 = ((~g21771));
assign g11511 = ((~II18509));
assign II15262 = ((~g481));
assign g13208 = ((~g9670));
assign g5944 = ((~g2151));
assign g12259 = ((~II19432));
assign g6080 = ((~II14587));
assign g26905 = ((~g26096)&(~g22319));
assign II38462 = ((~g29120));
assign g25573 = ((~II33396));
assign II27017 = ((~g19170));
assign g22615 = ((~g21900)&(~g18990));
assign g25198 = (g24691&g16651);
assign g13225 = ((~g9873));
assign g15800 = ((~g12909));
assign g23547 = (g8062&g22405);
assign g5749 = ((~II14195));
assign II28959 = ((~g21636));
assign g23611 = (g6194&g22509);
assign g20020 = (g18109&g18024&II26464);
assign g12499 = ((~g9074)&(~g9090)&(~g9101));
assign II38620 = ((~g29246));
assign II21301 = ((~g12438));
assign II40874 = ((~g30751));
assign g29422 = ((~II38647));
assign II32668 = ((~g18247))|((~g23999));
assign g18987 = ((~g15794));
assign g8791 = ((~II15989));
assign g8271 = ((~II15481));
assign g21890 = ((~g13530)&(~g19307));
assign g23368 = ((~g23135))|((~g22288));
assign g13144 = ((~g9968))|((~g7426));
assign g7643 = ((~g316));
assign g20371 = ((~g17471));
assign g27806 = ((~II36267));
assign II15902 = ((~g6486));
assign g27896 = ((~g27632)&(~g1222));
assign g21172 = (g19389&g19368&II27733);
assign II23874 = ((~g15797));
assign II22687 = ((~g14650));
assign II36668 = ((~g14966))|((~II36666));
assign g22793 = (g14472&g21647);
assign g21193 = (g20120&g16599&g16554);
assign II39761 = ((~g30072));
assign II15853 = ((~g3494));
assign II16814 = ((~g6486));
assign g10312 = (g5512&g4688);
assign g5884 = (g2400&g2469);
assign g29774 = ((~g29475)&(~g29211));
assign g25370 = ((~g24820));
assign g28684 = ((~II37599));
assign g27987 = ((~II36462));
assign II26237 = ((~g16857));
assign g10157 = (g7015&g4406);
assign g6087 = ((~g1186));
assign g5423 = ((~g2879));
assign II38412 = ((~g28720));
assign g27555 = ((~II35957));
assign g26363 = (g4894&g25643);
assign g27255 = ((~g26969)&(~g26233));
assign g12536 = ((~g8678));
assign g22114 = ((~g21372)&(~g19672));
assign g16969 = (g7888&g15220);
assign g16718 = ((~g14773)&(~g12531));
assign g20396 = ((~II26819));
assign g20964 = ((~g19760)&(~g17716));
assign II20595 = ((~g13271));
assign II36144 = ((~g27548));
assign II34656 = ((~g26173));
assign g19483 = ((~g16758));
assign II24538 = ((~g14268))|((~II24537));
assign g26792 = ((~g26451))|((~g3774));
assign II36459 = ((~g27258));
assign II31535 = ((~g23730));
assign g8964 = ((~II16270));
assign g17265 = ((~II23351));
assign g20659 = ((~II27250));
assign g16523 = ((~g14273));
assign g16099 = ((~g12844));
assign g6036 = ((~g2267));
assign g19103 = ((~g18590))|((~g2924));
assign g11666 = ((~g9098)&(~g9106)&(~g9113));
assign g29669 = ((~g29528)&(~g29300));
assign g12161 = ((~g8360));
assign g23268 = ((~II30257));
assign g22171 = ((~g21454)&(~g19789));
assign g10284 = (g6643&g4603);
assign g18823 = ((~g15182));
assign g21991 = ((~g21501))|((~g21536));
assign II29912 = ((~g23065));
assign II25671 = ((~g2160))|((~g18469));
assign g28430 = (g28128&g9196);
assign II31457 = ((~g23773));
assign II22860 = ((~g14885));
assign g24672 = (g24097)|(g20858);
assign g26248 = ((~II34198));
assign g23822 = (g14148&g23037);
assign g29344 = (g29076&g29065);
assign II17989 = ((~g3254));
assign g29717 = ((~g29583)&(~g1910));
assign g29286 = ((~g28807));
assign g24877 = ((~II32576))|((~II32577));
assign II14219 = ((~g801));
assign g28492 = (g18509&g28186);
assign g24657 = ((~g23723)&(~g22632));
assign g30508 = ((~II40104));
assign II13937 = ((~g1727));
assign g18308 = ((~g16174)&(~g6832));
assign g16551 = ((~g14395)&(~g14546));
assign II21137 = ((~g11749));
assign gbuf141 = (g1753);
assign g30102 = (g29849&g11348);
assign g30955 = ((~g30918)&(~g30945));
assign g15791 = ((~g12711))|((~g7085));
assign g7673 = ((~g319));
assign g26007 = ((~II33873));
assign II35443 = ((~g26757));
assign g29237 = ((~II38330));
assign g27608 = ((~g27152));
assign II33415 = ((~g24449));
assign g27239 = ((~II35554));
assign g21410 = (g6363&g20402);
assign g24047 = ((~g23023));
assign g22422 = ((~II28966));
assign g13489 = (g6026&g12219);
assign g28132 = ((~II36808));
assign II29135 = ((~g21804));
assign g19870 = (g686&g18927);
assign g13860 = (g7593&g12742);
assign II20589 = ((~g11629));
assign II32904 = ((~g24531));
assign g15222 = ((~II21505));
assign II27053 = ((~g19190));
assign II19415 = ((~g10549));
assign g20376 = ((~g16865)&(~g13787));
assign g7688 = ((~g1695));
assign g11520 = ((~II18536));
assign g22254 = (g21716&g12239);
assign g17965 = (g5009&g15582);
assign II40796 = ((~g30829));
assign g25193 = (g24653&g16626);
assign II32967 = ((~g25124));
assign g17249 = ((~II23335));
assign g22654 = (g21921&g12798);
assign g15900 = ((~g12711))|((~g6838));
assign g29646 = ((~II39056));
assign II16511 = ((~g6713));
assign II28189 = ((~g14079))|((~g19444));
assign g20132 = (g18593&g3182);
assign g7594 = ((~g2165));
assign g21623 = ((~II28152));
assign g8928 = ((~II16218));
assign II17042 = (g5976&g4860&g4861&g5334);
assign g5252 = ((~g1966));
assign g14690 = (g7841&g13101);
assign g4023 = ((~g702));
assign g17447 = (g4115&g15106);
assign II29978 = ((~g22670));
assign g28764 = ((~II37725));
assign II35416 = ((~g26884));
assign g16879 = (g15813&g8693);
assign II16123 = ((~g5406));
assign g27177 = ((~g26501));
assign g19235 = (g18478)|(g18611);
assign g19879 = (g2052&g18933);
assign g10531 = (g3806&g2647);
assign g30663 = ((~g16357)&(~g30472));
assign g24272 = ((~II31490));
assign g28428 = (g17825&g28155);
assign II28743 = ((~g13530))|((~II28741));
assign g28556 = (g27751)|(g25853);
assign II17765 = ((~g7976));
assign II37155 = ((~g28119));
assign g22509 = ((~II29055));
assign g17764 = ((~II23839));
assign g12894 = ((~g8934));
assign g25881 = (g2908&g25126);
assign g20113 = (g16836&g3142);
assign g25929 = ((~g24978))|((~g6713));
assign g15741 = ((~II21989));
assign g18635 = ((~II24744))|((~II24745));
assign g16054 = ((~g12783));
assign g15978 = ((~g11737)&(~g7152));
assign g29230 = ((~II38321));
assign g13149 = ((~g8676)&(~g8687)&(~g8703));
assign II32469 = ((~g17903))|((~II32468));
assign g24808 = ((~II32369))|((~II32370));
assign g29449 = ((~II38728));
assign g16781 = ((~g15003));
assign g21249 = ((~g19972));
assign g5869 = ((~g1615));
assign g8906 = (g7053&g1871);
assign g18849 = ((~g15311));
assign g6367 = ((~g285));
assign II37131 = ((~g28091));
assign g10772 = ((~g6978));
assign g21051 = ((~g19895)&(~g18088));
assign g5587 = ((~g3091));
assign II41011 = ((~g30775))|((~II41010));
assign g18478 = ((~II24513))|((~II24514));
assign g20469 = ((~II26910));
assign II20839 = ((~g13143));
assign II32400 = ((~g17927))|((~g24036));
assign II22604 = ((~g15080));
assign g19304 = ((~II25644))|((~II25645));
assign g25974 = ((~g24604)&(~g23527));
assign II23277 = ((~g9941))|((~g14320));
assign gbuf131 = (g1665);
assign g21764 = ((~g20228))|((~g6574));
assign g28390 = ((~II37319));
assign g28300 = ((~II37149));
assign g25623 = ((~II33448));
assign g28389 = (g2120&g27794);
assign g23636 = (g4191&g22537);
assign g29203 = (g15118&g28755);
assign II33583 = ((~g25068));
assign g27241 = (g10730&g26934);
assign g20139 = (g16836&g3151);
assign II21865 = ((~g13115));
assign II31121 = ((~g23017));
assign g27471 = ((~g23138)&(~g26764)&(~g24435));
assign g19242 = (g14244)|(g16501);
assign g24963 = ((~II32725))|((~II32726));
assign g22168 = ((~g21447)&(~g19781));
assign g25211 = ((~g24750)&(~g23558));
assign II15992 = ((~g6055));
assign II23047 = ((~g13894))|((~II23045));
assign g26670 = ((~g25362)&(~g17166));
assign g11004 = ((~II17913));
assign II29559 = ((~g21034));
assign g30400 = ((~g29997)&(~g30127));
assign g5648 = ((~II14104));
assign g8752 = ((~II15942));
assign II40994 = ((~g30795));
assign g25450 = ((~g16018)&(~g25086));
assign g30275 = ((~g16413)&(~g30109));
assign g17079 = (g8156&g15560);
assign g13328 = ((~g10334));
assign g9924 = (g6574&g4162);
assign g22258 = ((~g20679));
assign g23574 = ((~II30648));
assign II19667 = ((~g10822));
assign g25997 = ((~II33843));
assign g26466 = ((~II34428));
assign II31188 = ((~g21989));
assign II36873 = ((~g27971));
assign g10892 = ((~II17765));
assign II38226 = ((~g29108));
assign II16504 = ((~g3306));
assign g18784 = ((~g15037));
assign g11556 = ((~II18644));
assign g17396 = (g4020&g15037);
assign g21369 = (g15188&g20368);
assign II23056 = ((~g9264))|((~II23055));
assign g20362 = ((~g17433));
assign g18012 = (g5061&g15609);
assign II21461 = ((~g13052));
assign g12607 = ((~II19753));
assign II38832 = ((~g29324))|((~II38831));
assign g22871 = ((~II29669));
assign II40016 = ((~g30251));
assign g6677 = ((~II14808));
assign g29442 = ((~II38707));
assign g7476 = ((~g785));
assign g4389 = ((~g1512));
assign II15995 = ((~g7577));
assign gbuf81 = (g969);
assign g5369 = ((~g1423));
assign II14357 = ((~g785));
assign II20486 = ((~g10889));
assign g14910 = ((~g12207));
assign g4735 = ((~II13601));
assign II35992 = ((~g27106))|((~g15074));
assign g24070 = ((~g22812))|((~g14011));
assign II19803 = ((~g10754));
assign g29069 = ((~II38028));
assign II38869 = ((~g29181));
assign g19356 = (g18063&g3112);
assign II40194 = ((~g30370));
assign g9003 = ((~II16321));
assign g10382 = (g7162&g4791);
assign g27531 = ((~g26760)&(~g25181));
assign g17698 = ((~II23782));
assign g5615 = ((~II14073));
assign g21626 = (g13983&g14390&g19876&II28155);
assign II28509 = ((~g21427));
assign II14446 = ((~g3230));
assign g28494 = (g18474&g28018);
assign II31883 = ((~g23767));
assign II40934 = ((~g30827));
assign g29620 = ((~g14039)&(~g29262));
assign g7736 = ((~g1698));
assign g26547 = ((~g13796)&(~g25278));
assign g7479 = ((~g1861));
assign g12837 = ((~II19898));
assign g11699 = ((~g9822))|((~g3678));
assign g8614 = ((~II15800));
assign g3244 = ((~II13128));
assign g24151 = ((~g22530));
assign II23403 = ((~g13478));
assign g11141 = ((~II18055));
assign g4791 = ((~g1401));
assign g21367 = (g9203&g20366);
assign g21291 = (g9293&g20279);
assign g25684 = ((~g25106)&(~g6216));
assign II22797 = ((~g14165));
assign g9293 = ((~g5703));
assign g17144 = (g7958&g15724);
assign g16004 = (g5587&g11734);
assign g12115 = ((~g11462));
assign II24029 = ((~g6201))|((~II24028));
assign g26397 = (g5030&g25703);
assign II17933 = ((~g3254));
assign g7799 = ((~g1704));
assign g30443 = ((~II39997));
assign g22068 = ((~g21336)&(~g19606));
assign g9242 = ((~II16504));
assign g5877 = ((~g2294));
assign g19574 = (g8191&g17304);
assign g3306 = ((~II13165));
assign g16490 = ((~II22572));
assign II41018 = ((~g30768))|((~II41017));
assign g27985 = (g14342&g27489);
assign g29961 = (g29776&g29057);
assign g21238 = ((~g19954)&(~g5890));
assign g21502 = ((~g20525)&(~g16445));
assign II16041 = ((~g6486));
assign g22866 = ((~II29660));
assign II38924 = ((~g29205));
assign g25323 = ((~g24920));
assign II16569 = ((~g6000));
assign g30862 = ((~II40838));
assign II35716 = ((~g26865))|((~II35714));
assign g29681 = ((~g29555)&(~g29332));
assign g14483 = ((~g12170));
assign g25223 = ((~g24769)&(~g23579));
assign g22651 = ((~g21912)&(~g18997));
assign II20033 = ((~g9883))|((~II20031));
assign II26455 = (g18424)|(g18346)|(g18270);
assign g30258 = ((~g16291)&(~g30092));
assign g19799 = (g17640&g18074&II26240);
assign g10538 = (g7426&g5129);
assign g9631 = (g6314&g3925);
assign g16992 = ((~II22937))|((~II22938));
assign II35031 = ((~g26529));
assign g22358 = (g21782&g12389);
assign g11936 = ((~g11213));
assign II36627 = ((~g27302));
assign g11568 = ((~II18680));
assign g15837 = ((~g12657))|((~g6783));
assign g30397 = (g30241&g9019);
assign g22128 = ((~g21391)&(~g19703));
assign g29339 = ((~II38524));
assign g5962 = ((~g957));
assign g23518 = ((~g22914))|((~g14584))|((~g10735));
assign g13654 = (g8093&g11791);
assign g30575 = ((~g30412));
assign g28277 = ((~II37080));
assign g5790 = ((~g2129));
assign II39130 = ((~g29580));
assign II25971 = ((~g16671));
assign g21070 = ((~g19920)&(~g18204));
assign g22211 = (g21661&g12027);
assign g23299 = ((~II30350));
assign II35698 = ((~g26897));
assign g21160 = (g20120&g14478);
assign g13199 = ((~g9588));
assign g13046 = ((~g10814));
assign g22845 = ((~g19441))|((~g20885));
assign g23000 = ((~g16909)&(~g21067));
assign g5963 = ((~g1462));
assign g12943 = ((~g8984));
assign g28022 = ((~II36533));
assign II27593 = ((~g20025));
assign II33843 = ((~g25724));
assign II29288 = ((~g20939));
assign g29219 = ((~g28948)&(~g28474));
assign g22583 = ((~II29145));
assign g30112 = (g29861&g11432);
assign g17773 = (g4693&g15426);
assign II35455 = ((~g26881));
assign II17807 = ((~g8107));
assign g22221 = ((~g21932));
assign II17860 = ((~g5765));
assign g23386 = ((~g22483)&(~g21388));
assign II32576 = ((~g18155))|((~II32575));
assign g21324 = (g9391&g20323);
assign g30793 = ((~II40637));
assign II37815 = ((~g28391))|((~II37813));
assign g18893 = ((~g15467));
assign g15879 = ((~g12565))|((~g6232));
assign g15714 = ((~II21962));
assign g17482 = ((~II23570));
assign g21611 = (g7471&g19915);
assign g26781 = ((~g26044)&(~g10133));
assign II35756 = ((~g27117));
assign g7530 = ((~g496));
assign g26313 = ((~g25324));
assign g26236 = (g25899&g9371);
assign II17951 = ((~g6519));
assign g5730 = (g1012&g1066);
assign g8386 = (g6314&g234);
assign II24427 = ((~g7134))|((~II24426));
assign g14119 = ((~g11955));
assign g8120 = ((~g3197));
assign g12194 = ((~g10434)&(~g10494)&(~g10556));
assign g27480 = ((~II35824));
assign g23803 = ((~II31031));
assign g22494 = ((~II29040));
assign g12153 = ((~g10380)&(~g10445)&(~g10509));
assign II24575 = ((~g6216))|((~g14614));
assign gbuf103 = (g1209);
assign g30556 = ((~II40248));
assign g27842 = ((~g27632)&(~g1217));
assign g21935 = ((~II28450));
assign II36066 = ((~g27479));
assign II24149 = ((~g7079))|((~II24148));
assign g17476 = ((~II23564));
assign II30486 = ((~g23022));
assign g5862 = ((~g936));
assign g25127 = ((~g23525)&(~g22363));
assign II15239 = ((~g2966))|((~II15237));
assign g15903 = ((~g13404))|((~g12392));
assign II40534 = ((~g30693));
assign g24402 = ((~II31880));
assign g13257 = ((~II20310));
assign g21251 = (g19681&g15003&g16743);
assign II38428 = ((~g28732));
assign gbuf115 = (g1235);
assign II30392 = ((~g22226));
assign g12553 = ((~g8708));
assign g23907 = (g18436&g23079);
assign II38848 = ((~g29167));
assign g26648 = ((~g25821));
assign g17372 = ((~II23460));
assign g10672 = (g7391&g2682);
assign II37508 = ((~g27769));
assign g19789 = (g4561&g17701);
assign g23143 = ((~g21825));
assign II29122 = ((~g20742));
assign g30438 = (g30147&g11085);
assign g27101 = (g22157&g26654);
assign g25520 = (g24813)|(g23145);
assign g5795 = ((~g2376));
assign g10690 = (g3806&g2685);
assign g24916 = ((~g23502));
assign II30617 = ((~g22032));
assign II17705 = ((~g6836));
assign g28417 = ((~g24712)&(~g27830));
assign g30873 = ((~II40871));
assign II18341 = ((~g5610));
assign g24855 = (g18174&g23731);
assign II35518 = ((~g26959));
assign g29412 = ((~II38617));
assign g11951 = ((~g11240));
assign g9626 = ((~II16723));
assign g27204 = ((~II35449));
assign g17701 = ((~II23785));
assign g5701 = ((~II14149));
assign g9019 = ((~II16341));
assign g24712 = (g13585&g24153);
assign g29721 = ((~g6104)&(~g29583)&(~g25323));
assign g23681 = (g4310&g22573);
assign II31607 = ((~g23595));
assign g28218 = ((~II36903));
assign II29439 = ((~g20993));
assign II32868 = ((~g25118));
assign g8169 = ((~g2947));
assign II39794 = ((~g30130));
assign g15595 = (g5149&g13250);
assign g4711 = ((~g2235));
assign II36153 = ((~g27562));
assign g18630 = ((~g14483)&(~g16171));
assign g8888 = ((~II16156));
assign g25735 = ((~II33564));
assign g16127 = (g1678&g11813);
assign g30474 = ((~II40044));
assign II28126 = (g13963&g14360&g14016);
assign g16540 = ((~II22618));
assign g27993 = ((~II36476));
assign g28034 = ((~II36563));
assign g15513 = ((~II21772));
assign g28667 = (g27964&g13852);
assign II29386 = ((~g20973));
assign g30905 = ((~II40967));
assign g10256 = (g3722&g4561);
assign g16923 = (g7352&g15048);
assign g22708 = ((~g16113))|((~g21278));
assign g18808 = ((~g15115));
assign g19587 = (g8212&g17318);
assign g29671 = ((~g29534)&(~g29310));
assign g11725 = ((~g9968))|((~g3834));
assign g24094 = ((~g22339));
assign g23037 = ((~g21561));
assign g26342 = (g4818&g25606);
assign g5635 = ((~g2170));
assign g19633 = (g1319&g18809);
assign g21077 = (g20223&g12094);
assign g17315 = ((~II23403));
assign g30978 = ((~II41108));
assign g15981 = ((~g11687));
assign g24307 = ((~II31595));
assign g11659 = ((~II18845));
assign g6149 = ((~g3097));
assign g7545 = ((~g2920));
assign g20595 = ((~II27110));
assign g23469 = ((~II30511));
assign g8311 = ((~II15517));
assign g23124 = ((~g17129)&(~g21195));
assign g13579 = ((~II20799));
assign g28476 = (g26131&g28173);
assign g10228 = (g5512&g1810);
assign g30036 = ((~g29912));
assign g11577 = ((~II18707));
assign II29530 = ((~g21025));
assign g2636 = ((~II13098));
assign g30530 = ((~II40170));
assign g24750 = (g15454&g24104);
assign g24868 = ((~II32547))|((~II32548));
assign g16943 = ((~g13589));
assign g7558 = ((~g2165));
assign II15847 = ((~g3878));
assign g26973 = (g6301&g26226);
assign II21208 = ((~g11749));
assign g20189 = (g16825&g9289);
assign g29999 = (g29924&g22279);
assign g8463 = (g3254&g246);
assign g15998 = (g5469&g11732);
assign g15104 = (g4220&g13167);
assign g23318 = ((~II30407));
assign g5739 = (g1712&g1732);
assign g16029 = (g12071&g10877);
assign II25371 = ((~g18719));
assign g11534 = ((~II18578));
assign g8948 = ((~II16252));
assign g9811 = (g6574&g4070);
assign g24434 = ((~g23401)&(~g10238));
assign g21388 = (g6201&g19657);
assign g27306 = ((~g27046)&(~g26384));
assign g18964 = ((~g15741));
assign II22737 = ((~g14630));
assign gbuf168 = (g2006);
assign g28029 = ((~g26033)&(~g27247));
assign g26032 = (g25379&g19415);
assign g7557 = ((~g1874));
assign II36476 = ((~g27263));
assign g23620 = ((~II30738));
assign II23751 = ((~g14966));
assign g27109 = (g22157&g26658);
assign g20949 = ((~g19741)&(~g17673));
assign g14385 = ((~g12970));
assign g24352 = ((~II31730));
assign g30091 = (g29844&g11202);
assign II22745 = ((~g14725));
assign g4231 = ((~g708));
assign g16543 = ((~g14347));
assign II39258 = ((~g29696));
assign g22940 = ((~g19512))|((~g20956));
assign g8571 = ((~g3710))|((~g3678));
assign g25042 = ((~g24234)&(~g17031));
assign g19302 = ((~g17025));
assign g25299 = (g5659&g24850);
assign II33717 = ((~g24548));
assign g5941 = ((~g1639));
assign g10315 = (g7053&g1949);
assign g26281 = ((~II34241));
assign g19036 = ((~II25171));
assign II14298 = ((~g3217));
assign g11561 = ((~II18659));
assign g22758 = ((~II29496));
assign g18330 = (g5323&g15774);
assign g8464 = (g6314&g252);
assign g11975 = ((~g10107)&(~g10197)&(~g10282));
assign g30379 = ((~II39942));
assign g10789 = ((~g5650)&(~g5677)&(~g5709));
assign g5986 = ((~g960));
assign g5666 = ((~g216));
assign II16289 = ((~g5421));
assign II20700 = ((~g12450));
assign II13236 = ((~g2703));
assign g30410 = (g30139&g11028);
assign II28913 = ((~g21255));
assign II39573 = ((~g29936));
assign II33903 = ((~g25880));
assign g22073 = ((~g21337)&(~g19616));
assign g4696 = ((~g2089));
assign g23887 = ((~g22328));
assign g24227 = ((~g22270)&(~g21137));
assign g26865 = ((~II35035))|((~II35036));
assign g27284 = ((~g27018)&(~g26334));
assign II25180 = ((~g18992));
assign g18536 = ((~g14520));
assign g29568 = ((~II38958));
assign g24374 = ((~II31796));
assign g8530 = ((~g6156));
assign g21961 = ((~II28509));
assign g28370 = ((~II37269));
assign g11860 = ((~g9765)&(~g9893)&(~g10012));
assign gbuf6 = (g2818);
assign g19505 = ((~g16895));
assign II33390 = ((~g25038));
assign g20850 = ((~g19468));
assign II28273 = ((~g19515))|((~II28271));
assign g6054 = ((~II14541));
assign g27726 = (g27531&g20732);
assign II16961 = ((~g7303));
assign g22716 = ((~II29402));
assign g23462 = (g17988&g22609);
assign g10200 = (g6486&g587);
assign g7694 = ((~g1784));
assign II20670 = ((~g12552));
assign g12134 = ((~g8321));
assign g9126 = (g3774&g7779);
assign g21087 = ((~II27646));
assign g24346 = ((~II31712));
assign g27137 = ((~g26202));
assign g28360 = ((~g15725)&(~g28098));
assign g26278 = (g4541&g25515);
assign II16465 = ((~g6000));
assign II30281 = ((~g22635));
assign g19773 = (g1339&g17670);
assign g20923 = ((~g19699)&(~g17578));
assign g11587 = ((~II18737));
assign g26915 = ((~g25708))|((~g26327))|((~g25648));
assign g14124 = ((~g12899));
assign II25533 = ((~g52))|((~II25532));
assign g28623 = ((~g27872));
assign II15590 = ((~g3410));
assign II32334 = ((~g18131))|((~II32333));
assign g9640 = ((~II16741));
assign g28401 = (g7782&g27831);
assign II16827 = (g5771&g5987&g4911&g4912);
assign g20583 = ((~II27074));
assign g23608 = ((~II30716));
assign g27723 = (g27464&g20679);
assign g22639 = ((~II29243));
assign g26723 = ((~II34776));
assign g24767 = (g15540&g24121);
assign g21643 = ((~g16591)&(~g19987));
assign g29819 = (g29751&g22294);
assign g29365 = ((~g28900));
assign g9941 = ((~g6035));
assign II36267 = ((~g27395));
assign g13649 = ((~g11711));
assign g12071 = ((~g10783));
assign g22731 = ((~II29435));
assign g4876 = ((~g2785));
assign II18223 = ((~g6448));
assign g25189 = ((~g24502)&(~g10133));
assign g11746 = ((~g10895));
assign g29800 = ((~II39252));
assign g21080 = ((~g19935)&(~g18311));
assign g9815 = ((~g5598));
assign g24030 = ((~II31250));
assign II21310 = ((~g12332));
assign g5089 = ((~g2093));
assign g17291 = ((~II23377));
assign g27379 = ((~II35702))|((~II35703));
assign g24636 = ((~g24183)&(~g530));
assign g12207 = ((~g10443)&(~g10507)&(~g10566));
assign g19265 = ((~g16572));
assign g27587 = ((~g26897))|((~g2124));
assign g17382 = (g8252&g16002);
assign g17233 = ((~II23317));
assign g24423 = ((~II31943));
assign g4323 = ((~II13421));
assign gbuf16 = (g2848);
assign II22554 = ((~g14765));
assign II15983 = ((~g3878));
assign g18061 = (g5138&g15652);
assign g24801 = ((~II32356))|((~II32357));
assign g19624 = (g4003&g17387);
assign g27274 = ((~g27002)&(~g26309));
assign g20915 = ((~g19674)&(~g17542));
assign g27552 = (g23974&g27162);
assign II17954 = ((~g6369));
assign g18584 = ((~g16230)&(~g14570));
assign II40838 = ((~g30822));
assign g8473 = (g6783&g1615);
assign II40510 = ((~g30686));
assign g13750 = ((~g12439));
assign g27440 = ((~II35780));
assign II34665 = ((~g26191));
assign g30613 = ((~g30412)&(~g2607));
assign g10934 = ((~II17825));
assign g4318 = ((~g2800));
assign g19084 = ((~g16586))|((~g16602));
assign g6836 = ((~g1666));
assign II22938 = ((~g13906))|((~II22936));
assign g24866 = ((~II32539))|((~II32540));
assign II24689 = (g14811&g14910&g16201);
assign g17509 = (g4228&g15182);
assign g10299 = (g6713&g1128);
assign g12158 = ((~g8351));
assign g18105 = ((~g14719));
assign g26965 = (g23320&g26540);
assign g25851 = ((~II33695));
assign g15185 = ((~II21482));
assign g25982 = ((~II33798));
assign g23590 = (g4009&g22477);
assign g30307 = ((~II39764));
assign II36885 = ((~g28003));
assign g9159 = ((~II16457));
assign g21424 = (g9277&g20415);
assign g5853 = ((~g246));
assign g29506 = ((~II38848));
assign II30776 = ((~g22079));
assign g19276 = ((~II25572))|((~II25573));
assign II25041 = ((~g14895));
assign g30139 = ((~g30011));
assign g12066 = ((~g11404));
assign g29384 = ((~g29002));
assign g15237 = ((~II21520));
assign II23113 = ((~g9356))|((~g13848));
assign g12762 = ((~II19826));
assign g10513 = (g6980&g5064);
assign g26439 = ((~II34400));
assign g30842 = ((~II40778));
assign g29977 = ((~II39469));
assign II13974 = ((~g1769));
assign g9079 = (g5473&g7655);
assign g27019 = (g23364&g26587);
assign g25206 = ((~g24746)&(~g23550));
assign II30483 = ((~g23126));
assign g29271 = ((~g28764));
assign g27055 = (g22005&g26621);
assign g20916 = ((~g19675)&(~g17543));
assign g24469 = ((~g23955))|((~g3494));
assign g11623 = ((~g10961));
assign II14519 = ((~g1158));
assign g22020 = (g2366&g21225);
assign g11705 = ((~g9968))|((~g3834));
assign g11570 = ((~II18686));
assign g9137 = (g7015&g7799);
assign g23067 = ((~g17015)&(~g21122));
assign g28489 = ((~g26756)&(~g27720));
assign g22749 = ((~II29481));
assign g27918 = ((~II36379));
assign g12333 = ((~II19500));
assign g9778 = (g6369&g4035);
assign II34411 = ((~g25268));
assign g14958 = (g4016&g13153);
assign g28914 = (g14092&g28643);
assign g29405 = ((~II38602));
assign g24311 = ((~II31607));
assign II20709 = ((~g13070));
assign II21830 = ((~g13129));
assign g30368 = ((~II39913));
assign g18870 = ((~g15393));
assign II28476 = ((~g21064));
assign II17972 = ((~g7558));
assign II32916 = ((~g24597));
assign II32431 = ((~g17815))|((~II32430));
assign g11895 = ((~g11144));
assign g15207 = ((~II21497));
assign g11772 = ((~g9383)&(~g9462)&(~g9580));
assign II24436 = ((~g14153))|((~g15022));
assign g27621 = ((~g27188)&(~g17100));
assign g12829 = ((~g8874));
assign g24417 = ((~II31925));
assign g30116 = (g29921&g22236);
assign g25973 = (g24847&g13838);
assign g19349 = ((~g16647));
assign g12769 = ((~II19833));
assign g20893 = ((~g19628)&(~g17449));
assign g18037 = (g5095&g15631);
assign g15572 = (g4973&g12860);
assign II36327 = ((~g27413));
assign g7578 = ((~g1846));
assign II30959 = ((~g22138));
assign g23092 = ((~g17055)&(~g21154));
assign g4201 = ((~g2851));
assign g4535 = ((~g1541));
assign g16341 = ((~g12377))|((~g12407));
assign g27767 = ((~g27561)&(~g27107));
assign g29231 = ((~g29022)&(~g28494));
assign g9522 = (g6314&g8203);
assign g4088 = ((~II13316));
assign g24694 = ((~g24183)&(~g534));
assign g23493 = ((~g22203));
assign g13466 = ((~II20697));
assign g30522 = ((~II40146));
assign g26432 = (g5145&g25767);
assign g30867 = ((~II40853));
assign II32203 = ((~g23528));
assign g17118 = ((~g13915))|((~g13893));
assign g29208 = (g15188&g28764);
assign g13439 = ((~II20616));
assign g8474 = (g6574&g1621);
assign g16094 = ((~g6631)&(~g12499)&(~g10952));
assign II25105 = ((~g18959));
assign g29533 = (g28762&g29373);
assign II26025 = ((~g16803));
assign g25961 = (g24770&g11901);
assign g26027 = (g25418&g22271);
assign g22059 = ((~g21324)&(~g19591));
assign II33564 = ((~g24461));
assign g23302 = ((~II30359));
assign g16161 = (g1202&g11837);
assign g5688 = (g1012&g1051);
assign g28909 = (g14062&g28642);
assign g13057 = ((~g10784));
assign g24291 = ((~II31547));
assign g25484 = ((~II33312));
assign II39077 = ((~g29563));
assign II24038 = ((~g9374))|((~II24036));
assign g16135 = (g12187&g10980);
assign g29194 = ((~g14958)&(~g28881));
assign II22120 = ((~g12909));
assign g10707 = (g7162&g5355);
assign II33630 = ((~g25071));
assign g26591 = ((~g25612));
assign g26533 = ((~g25454));
assign g8893 = ((~II16163));
assign II20334 = ((~g9067));
assign g28085 = ((~II36696));
assign II27191 = ((~g20470));
assign g20799 = ((~II27388));
assign g3241 = ((~II13119));
assign g25764 = ((~g25076)&(~g21615));
assign g16049 = (g6638&g11763);
assign g17203 = ((~g13568));
assign g27223 = ((~II35506));
assign g28246 = ((~II36987));
assign g29076 = ((~g9391))|((~g28567));
assign g24792 = (g15694&g24143);
assign g15483 = ((~II21742));
assign g22609 = ((~g21108));
assign g30573 = ((~g30405));
assign g29988 = (g29881&g8382);
assign g25824 = ((~II33662));
assign g18883 = ((~g13846)&(~g12128));
assign g15993 = ((~g12926))|((~g7162));
assign g28084 = ((~II36693));
assign g18554 = ((~g13573));
assign II18485 = ((~g8809));
assign g22536 = ((~g17076)&(~g21911));
assign g20424 = ((~g17661));
assign II20048 = ((~g10185))|((~g10095));
assign gbuf194 = (g2470);
assign II16644 = ((~g5473));
assign g11548 = ((~II18620));
assign g25313 = ((~g24868));
assign II25722 = ((~g74))|((~II25721));
assign g27353 = ((~II35667));
assign g11969 = ((~g11268));
assign g8079 = ((~g1868));
assign II26630 = (g18744&g15080&g13774);
assign g28835 = ((~II37800));
assign g28931 = (g14153&g28645);
assign g9461 = (g3410&g8138);
assign g24467 = ((~g23803))|((~g3774));
assign g29541 = (g29214&g29379);
assign g24268 = ((~II31478));
assign g20008 = ((~g18977)&(~g7338));
assign g17369 = ((~II23457));
assign g6046 = ((~II14525));
assign II27705 = ((~g20545));
assign II34879 = ((~g26240));
assign g20499 = (g17648&g11933);
assign g21139 = (g19505)|(g16546)|(g14186);
assign g23764 = ((~II30953))|((~II30954));
assign g12968 = ((~g8520)&(~g8535)&(~g8548));
assign g20147 = (g16254&g13756&II26593);
assign g20504 = ((~g18355));
assign g21815 = (g18717)|(g20293)|(g20283)|(g18654);
assign II28318 = (g19092)|(g19088)|(g19079);
assign g20067 = ((~II26505));
assign g8617 = ((~II15803));
assign g16286 = (g5639&g13280);
assign g19419 = ((~II25856))|((~II25857));
assign g8008 = ((~g1168));
assign g5419 = ((~II13971));
assign g30787 = ((~g30594)&(~g22387));
assign g18864 = ((~g15382));
assign g10221 = (g6783&g4529);
assign g13789 = (g7140&g12554);
assign g28708 = (g28392&g22260);
assign g28638 = ((~g28200));
assign g11840 = ((~g9726)&(~g9810)&(~g9925));
assign II15448 = ((~g3237));
assign g29728 = ((~g6104)&(~g29583)&(~g25401));
assign gbuf88 = (g1039);
assign g27087 = (g22021&g26644);
assign g21885 = ((~g18556))|((~g19279))|((~g19297));
assign g26299 = (g4644&g25543);
assign g26016 = ((~II33900));
assign g26643 = ((~g25802));
assign g24318 = ((~II31628));
assign g6781 = ((~g970));
assign g19215 = (g18606)|(g18231);
assign g14657 = ((~II21252));
assign II16255 = ((~g3900));
assign g30709 = ((~g14228)&(~g30397));
assign gbuf69 = (g623);
assign g23831 = (g22962&g9673);
assign II41038 = ((~g30798));
assign g29374 = ((~g28951));
assign g25507 = ((~II33335));
assign g21756 = ((~g19070)&(~g18584));
assign gbuf90 = (g1052);
assign g7880 = ((~g3201));
assign II25915 = ((~g18025))|((~II25913));
assign g25435 = ((~II33257));
assign g4891 = ((~g583));
assign g11622 = ((~g8183)&(~g11332)&(~g7928)&(~g11069));
assign II19426 = ((~g10574));
assign gbuf13 = (g2839);
assign II38024 = ((~g28556));
assign II30695 = ((~g22056));
assign II41126 = ((~g30972));
assign g23644 = ((~II30786));
assign II25031 = ((~g8029))|((~II25030));
assign II35461 = ((~g26895));
assign g11839 = ((~g9724)&(~g9807)&(~g9922));
assign g14811 = ((~g12097));
assign g30567 = ((~g30403));
assign g23078 = ((~II29827));
assign g27080 = (g23377&g26637);
assign II30692 = ((~g22055));
assign g28127 = (g27622&g10409);
assign g30313 = ((~II39782));
assign II26898 = ((~g17248));
assign g29417 = ((~II38632));
assign g21771 = ((~g20255))|((~g6838));
assign g10572 = (g3618&g5170);
assign g13060 = ((~g10801));
assign g30700 = ((~g13952)&(~g30388));
assign II40008 = ((~g30250));
assign g25741 = ((~II33570));
assign g26052 = (g25941&g21087);
assign II30997 = ((~g22148));
assign g30516 = ((~II40128));
assign g23937 = ((~g22812))|((~g13918));
assign g5905 = ((~g1457));
assign g22771 = ((~g16223))|((~g21293));
assign g12327 = ((~g10639)&(~g10671)&(~g10689));
assign g29323 = (g29068&g28983);
assign g30910 = ((~II40982));
assign g24592 = ((~II32164));
assign g7727 = ((~g2390));
assign g23722 = (g4433&g22603);
assign g16454 = (g5990&g12158);
assign g30218 = (g30040&g8961);
assign g20104 = (g5391&g18619);
assign g22476 = ((~g21057));
assign g11481 = ((~g4204));
assign g26512 = ((~g25853));
assign II35087 = ((~g26667));
assign g22667 = (g14062&g21530);
assign II32146 = ((~g24219));
assign g15438 = ((~g12296));
assign g20302 = ((~g17282));
assign g18924 = ((~g15585));
assign g12407 = (g7573)|(g10779);
assign g24161 = ((~g22543));
assign g25259 = ((~g24853)&(~g23768));
assign g26554 = ((~g25502));
assign g7152 = ((~g3136));
assign g20719 = ((~II27308));
assign g15930 = ((~g12711))|((~g7085));
assign II21711 = ((~g13108));
assign II35741 = ((~g27118));
assign g19044 = ((~II25195));
assign g23606 = (g4070&g22500);
assign II28928 = ((~g21263));
assign II24493 = ((~g6301))|((~g14048));
assign II36444 = ((~g27482));
assign II24380 = ((~g6212))|((~g13978));
assign II26590 = (g14811&g18699&g18758);
assign II30260 = ((~g22743));
assign g12058 = ((~g11392));
assign g13453 = ((~II20658));
assign g21706 = ((~g20124)&(~g14431)&(~g14514));
assign II18623 = ((~g11003));
assign II37322 = ((~g27865))|((~g27855));
assign g25652 = ((~II33476));
assign g24102 = ((~g22418));
assign g15753 = (g7542&g12962);
assign II37656 = ((~g28365));
assign II23808 = ((~g9150))|((~II23806));
assign II38734 = ((~g29335));
assign g29524 = (g28739&g29365);
assign g23576 = ((~II30654));
assign g11478 = ((~II18444));
assign g11157 = ((~II18073));
assign g18933 = ((~g15625));
assign g4659 = ((~g1398));
assign g10303 = (g3522&g4656);
assign g20354 = ((~g17419));
assign g11468 = ((~II18432));
assign II38157 = ((~g28882));
assign g10994 = ((~II17895));
assign g8625 = (g3494&g7158);
assign g19714 = (g2020&g18844);
assign g5997 = ((~g2330));
assign g21400 = ((~g19918));
assign II19972 = (g9310&g9248&g9203&g9174);
assign g16481 = ((~II22545));
assign g23255 = ((~II30218));
assign g20287 = ((~g17252));
assign II39628 = ((~g30078));
assign II19787 = ((~g8726));
assign g9663 = (g3410&g3957);
assign g13150 = ((~g8287))|((~g3462));
assign II15887 = ((~g5693));
assign g19257 = (g18531)|(g18578);
assign g17892 = ((~g13954));
assign g14068 = ((~II21064));
assign g12087 = ((~g11435));
assign g4652 = ((~g1262));
assign g23599 = (g4041&g22487);
assign g8769 = ((~II15961));
assign g16615 = (g15971)|(g14753);
assign g5753 = ((~g228));
assign g6026 = ((~g2270));
assign g21801 = (g19128)|(g19608)|(g16686);
assign II25138 = ((~g18960));
assign g14775 = ((~II21313));
assign g24339 = ((~II31691));
assign g8100 = ((~g3070));
assign g26843 = ((~II34990));
assign g16591 = ((~g15933)&(~g15913)&(~g15890));
assign g29647 = ((~II39059));
assign g5549 = ((~II14027));
assign II21443 = ((~g12923));
assign g30893 = ((~II40931));
assign g26624 = ((~g25720));
assign II16372 = ((~g3774));
assign g16402 = (g5947&g12064);
assign II18773 = ((~g10830));
assign g28673 = ((~II37566));
assign g21958 = ((~II28500));
assign g30920 = (g30787&g22298);
assign II19549 = ((~g10683));
assign II37638 = ((~g28395));
assign g14637 = ((~g12329));
assign g9761 = (g6232&g4006);
assign g28014 = ((~g27373));
assign g5235 = ((~g1134));
assign g6060 = ((~II14559));
assign II24532 = ((~g14355))|((~II24530));
assign g20140 = ((~g16830));
assign II36702 = ((~g27322));
assign II23960 = ((~g14171))|((~II23958));
assign II29969 = ((~g22640));
assign g19163 = ((~g17486)&(~g15244));
assign g13580 = ((~II20802));
assign g10600 = (g7488&g5230);
assign g26181 = ((~II34083));
assign g18130 = (g5193&g15688);
assign II36307 = ((~g27400));
assign II32380 = ((~g24027))|((~II32378));
assign g8961 = ((~II16267));
assign II28693 = ((~g21847));
assign g12118 = ((~g11472));
assign g23790 = (g22958&g9592);
assign g13283 = ((~g10176));
assign g5275 = ((~g2659));
assign g4495 = ((~g869));
assign II37077 = ((~g28101));
assign g15644 = ((~II21897));
assign g27210 = ((~II35467));
assign g8546 = (g3254&g210);
assign g20634 = ((~II27225));
assign II32370 = ((~g24012))|((~II32368));
assign II25560 = ((~g56))|((~g17724));
assign g20432 = ((~g17688));
assign g29981 = (g29869&g8330);
assign g20408 = ((~g17594));
assign g6194 = ((~g2746));
assign g15452 = (g7916&g12808);
assign II24546 = ((~g9649))|((~II24544));
assign II31613 = ((~g23596));
assign II21537 = ((~g13071));
assign g25025 = ((~g23748))|((~g7015));
assign g30736 = (g30584&g20669);
assign g15527 = (g5034&g13233);
assign II23578 = ((~g15879));
assign g21650 = (g16551&g19524&g14301);
assign g27224 = ((~II35509));
assign g5760 = ((~g744));
assign II31463 = ((~g23774));
assign g27563 = ((~g26922)&(~g24708));
assign g19380 = ((~g16656));
assign g7590 = ((~g1155));
assign g8218 = ((~g858));
assign g15612 = ((~II21868));
assign g13036 = ((~g10831));
assign II36111 = ((~g27505));
assign g8987 = ((~II16303));
assign g20714 = ((~II27303));
assign g28329 = (g27823&g20708);
assign g22760 = ((~II29500));
assign II22820 = ((~g14402));
assign II18356 = ((~g7085));
assign g30696 = (g30383&g10943);
assign g16393 = (g5941&g12053);
assign g6067 = ((~II14580));
assign g18058 = (g5123&g15641);
assign II38434 = ((~g28735));
assign II20497 = ((~g8579));
assign g15805 = ((~g12565))|((~g6232));
assign g22297 = ((~g20757));
assign g29452 = ((~II38737));
assign II24228 = ((~g14316))|((~II24226));
assign g10352 = (g7488&g4728);
assign g20401 = ((~g17570));
assign g18561 = ((~II24647))|((~II24648));
assign II27349 = ((~g19431));
assign II26432 = (g18277&g18189&g18090);
assign g12507 = ((~g10213)&(~g10300)&(~g10376));
assign g24383 = ((~II31823));
assign g25471 = ((~II33297));
assign g29893 = ((~g29685));
assign g21379 = (g9427&g20379);
assign g23305 = ((~II30368));
assign II16147 = ((~g3878));
assign II26745 = (g18772&g18796&g16325);
assign II15372 = ((~g3129));
assign g6626 = ((~g2020));
assign II23493 = ((~g15846));
assign g12262 = ((~g10519)&(~g10581)&(~g10623));
assign II15271 = ((~g1186));
assign g26148 = ((~g8305))|((~g14753))|((~g25445))|((~g25413));
assign g15717 = (g7924&g13285);
assign g24816 = ((~II32388));
assign g22357 = ((~g20816));
assign II29638 = ((~g21063));
assign g12036 = ((~g10205)&(~g10292)&(~g10370));
assign II37999 = ((~g28584));
assign g5555 = ((~II14037));
assign g28852 = (g27875&g28623);
assign g19894 = ((~II26340));
assign g12063 = ((~g11395));
assign g24134 = ((~g22396));
assign g21278 = ((~II27827));
assign g9471 = ((~g5820));
assign g11517 = ((~II18527));
assign g29001 = ((~g9161))|((~g28512));
assign II18518 = ((~g8893));
assign II25084 = ((~g14885));
assign g30318 = ((~II39797));
assign g23188 = ((~II30017));
assign II25459 = ((~g18867));
assign II36647 = ((~g27308));
assign g26336 = ((~g25981)&(~g13481));
assign II40326 = ((~g30356));
assign g20606 = ((~II27143));
assign g30548 = ((~II40224));
assign II30722 = ((~g22063));
assign II15538 = ((~g6369));
assign g28767 = ((~g28452)&(~g27945));
assign g14419 = (g7779&g13003);
assign II23351 = ((~g15788));
assign g13179 = ((~g9387));
assign II26624 = (g14863&g18789&g13724);
assign g22101 = ((~g21361)&(~g19654));
assign g12756 = ((~II19820));
assign II25201 = ((~g16843));
assign g28645 = ((~g27952));
assign II24943 = ((~g14811));
assign g24549 = ((~II32081));
assign g22014 = ((~II28564));
assign g15491 = (g4954&g13222);
assign g13316 = (g5675&g11210);
assign g24668 = ((~g23482));
assign II34851 = ((~g26354));
assign g22290 = ((~g20739));
assign g14176 = ((~g11981));
assign g24077 = ((~II31298));
assign II21511 = ((~g13064));
assign g11684 = ((~g9676))|((~g3522));
assign g22305 = (g21742&g12340);
assign g7605 = ((~g1849));
assign g15407 = (g4778&g13207);
assign g29102 = ((~II38097));
assign II25338 = ((~g17746));
assign g26194 = ((~II34108));
assign II24428 = ((~g14332))|((~II24426));
assign g30917 = (g12446&g30766);
assign g17191 = ((~g14703))|((~g14725));
assign g28093 = ((~II36714));
assign II18244 = ((~g5720));
assign g26482 = ((~g25357))|((~g753));
assign II37164 = ((~g28125));
assign g21682 = ((~II28210));
assign g17086 = ((~g14691)&(~g15913)&(~g14650));
assign g10387 = (g3566&g4806);
assign II33918 = ((~g25763));
assign g23250 = ((~II30203));
assign g16369 = (g5916&g12002);
assign II31622 = ((~g23620));
assign g5977 = ((~g2612));
assign g13634 = (g12776&g8617);
assign II19211 = ((~g10486));
assign II22946 = ((~g15188))|((~II22945));
assign g20014 = (g7615&g16749);
assign g21787 = (g19121)|(g19578)|(g16665);
assign g5718 = ((~g903));
assign g20443 = ((~g17749));
assign g19049 = ((~II25210));
assign II30131 = ((~g22864));
assign g27494 = ((~II35844));
assign II14688 = ((~g2599));
assign g8360 = ((~II15562));
assign g11355 = ((~II18311));
assign g5420 = ((~II13974));
assign g13527 = (g6047&g12325);
assign g12467 = ((~g9034)&(~g9056)&(~g9065));
assign g28233 = ((~II36948));
assign II32265 = ((~g17903))|((~g23936));
assign g18446 = ((~g13741));
assign g5349 = ((~g2877));
assign II29033 = ((~g21741));
assign II21995 = ((~g13146));
assign g15080 = ((~g12305));
assign g26582 = ((~g25585));
assign g14677 = ((~II21259));
assign g11450 = ((~II18414));
assign II15873 = ((~g5655));
assign g5727 = ((~g989));
assign g6643 = ((~II14802));
assign g11791 = ((~II18969));
assign II18238 = ((~g5593));
assign g16000 = ((~g12984))|((~g7488));
assign g22207 = (g21278&g16910);
assign g4629 = ((~g820));
assign g24215 = ((~g16993)&(~g22254));
assign g13589 = ((~II20813));
assign g12248 = ((~g10508)&(~g10567)&(~g10612));
assign g27658 = ((~g26851)&(~g26068));
assign II36650 = ((~g27309));
assign II33551 = ((~g24510));
assign g25186 = (g24969)|(g24916);
assign g11580 = ((~II18716));
assign g23191 = ((~II30026));
assign II38909 = ((~g29198));
assign II34201 = ((~g25246));
assign g17951 = ((~II23992));
assign g29787 = ((~g29487)&(~g29240));
assign g8725 = (g7391&g7912);
assign g17313 = ((~g16109));
assign g30588 = ((~g6119)&(~g30412)&(~g25353));
assign II15893 = ((~g3834));
assign g23897 = ((~II31165));
assign II25415 = ((~g18835));
assign g25367 = ((~g24676));
assign II21755 = ((~g11704));
assign g25466 = (g6222&g24827);
assign g17124 = ((~g14725)&(~g15942)&(~g14677));
assign g24348 = ((~II31718));
assign II28087 = ((~g19184));
assign g4833 = ((~g2087));
assign g5756 = ((~g304));
assign II37736 = ((~g28567));
assign g28791 = ((~II37752));
assign II25074 = ((~g14301));
assign g24214 = ((~g16990)&(~g22250));
assign g15782 = ((~g13332))|((~g12354));
assign g30199 = ((~g30026));
assign gbuf153 = (g1944);
assign g27111 = (g5309&g26490);
assign g22409 = ((~II28953));
assign g27719 = (g27496&g20649);
assign g9097 = (g3618&g7688);
assign II31742 = ((~g23629));
assign II17715 = ((~g8107));
assign g23015 = ((~g21514));
assign g25336 = ((~II33168));
assign g10150 = (g6574&g4389);
assign II20490 = ((~g9067));
assign g12472 = ((~g8617));
assign g24827 = ((~II32419));
assign g20255 = ((~II26679));
assign g24452 = ((~g23923))|((~g3338));
assign g14217 = ((~g11999));
assign g5990 = ((~g1645));
assign g8841 = (g6486&g490);
assign g30685 = ((~g29992)&(~g30000)&(~g30372));
assign g13883 = ((~g11656));
assign II38014 = ((~g28584));
assign g13602 = ((~g12326));
assign g9144 = (g2986)|(g5389);
assign g12389 = ((~II19549));
assign g27262 = ((~g26981)&(~g26268));
assign II30404 = ((~g22948));
assign g20295 = ((~II26714));
assign g18905 = ((~g15516));
assign II18049 = ((~g6314));
assign g14719 = ((~g12288));
assign g25078 = ((~g23419)&(~g22201));
assign g30655 = ((~g16300)&(~g30458));
assign II37587 = ((~g28552));
assign g22035 = ((~g21303)&(~g19562));
assign g18971 = ((~II25021));
assign g8684 = ((~II15882));
assign g10580 = (g3650&g5176);
assign g11990 = ((~II19174));
assign g26851 = (g5741&g26313);
assign g15818 = ((~g13024))|((~g12354));
assign g17121 = ((~II23124))|((~II23125));
assign g21003 = ((~g19820)&(~g15506));
assign II18441 = ((~g5837));
assign g20513 = ((~II26960));
assign g20326 = (g13805&g16404&II26745);
assign g4398 = ((~g1545));
assign II13742 = ((~g1501));
assign g12514 = (g7848&g9140);
assign g7838 = ((~g477));
assign g28263 = ((~II37038));
assign g22146 = ((~g21412)&(~g19737));
assign g16514 = ((~II22604));
assign g11596 = ((~II18764));
assign II34719 = ((~g26238));
assign g24505 = ((~g23771)&(~g19825));
assign g21218 = (g20212&g12421);
assign II36046 = ((~g26957));
assign g12296 = ((~II19466));
assign g11554 = ((~II18638));
assign g13619 = (g6162&g12466);
assign g12462 = ((~II19648));
assign gbuf70 = (g626);
assign g27217 = ((~II35488));
assign g13342 = ((~II20417));
assign g20048 = (g16749&g3127);
assign g19548 = (g16974&g16820&g14936);
assign g4182 = ((~g2223));
assign g30003 = (g29901&g8469);
assign g30066 = ((~g29816)&(~g13517));
assign g30078 = ((~II39577));
assign g30457 = (g30151&g11216);
assign g29379 = ((~g28975));
assign g29839 = (g29747&g20827);
assign g9335 = ((~II16556));
assign II21566 = ((~g13077));
assign g4000 = ((~g153));
assign II36906 = ((~g27989));
assign g27764 = ((~g27541)&(~g27095));
assign g27463 = ((~II35803));
assign g23439 = ((~II30470));
assign II25067 = ((~g14565));
assign g28386 = ((~II37304))|((~II37305));
assign g28710 = (g28403&g22262);
assign g25245 = ((~g24809)&(~g23636));
assign g11529 = ((~II18563));
assign II24486 = ((~g14541))|((~II24485));
assign II27125 = ((~g19652));
assign g13122 = ((~g9968))|((~g7488));
assign II32285 = ((~g17815))|((~II32284));
assign g10357 = ((~II17311));
assign II28766 = ((~g21901))|((~II28765));
assign g19819 = (g18038&g16092);
assign g26136 = ((~II34032));
assign g8968 = ((~II16276));
assign g10179 = ((~II17143));
assign g28666 = (g27980&g12106);
assign g22740 = ((~II29456));
assign II33614 = ((~g24521));
assign g30183 = ((~g30022));
assign II40739 = ((~g30661));
assign g20451 = ((~g17779));
assign g3774 = ((~II13228));
assign g15392 = (g4753&g13206);
assign g9907 = (g6369&g4133);
assign II18198 = ((~g7896))|((~II18197));
assign II39866 = ((~g30279));
assign II20673 = ((~g13397));
assign g25170 = ((~II32988));
assign g26199 = ((~g25961)&(~g13291));
assign II30020 = ((~g22519));
assign g15651 = (g5135&g12904);
assign II14525 = ((~g1852));
assign g26440 = ((~g16595))|((~g25190));
assign II25557 = ((~g18957));
assign II38659 = ((~g29322));
assign II25624 = ((~g1466))|((~II25623));
assign II38456 = ((~g28747));
assign II27838 = ((~g19936));
assign g4610 = ((~g596));
assign II27352 = ((~g19358));
assign g28996 = (g14414&g28653);
assign II18145 = ((~g6519));
assign II36803 = ((~g27348));
assign g29214 = ((~g28931)&(~g28469));
assign II17658 = ((~g6367));
assign g10195 = (g5438&g4471);
assign g19948 = ((~g17896));
assign g20999 = ((~g19816)&(~g17853));
assign II36280 = ((~g27390));
assign g27510 = ((~II35872));
assign g17676 = ((~II23760));
assign g18062 = (g7462&g15655);
assign II15469 = ((~g3244));
assign II40640 = ((~g30569));
assign II40637 = ((~g30570));
assign g30692 = ((~g13498)&(~g30361));
assign g10042 = (g3410&g4237);
assign II29067 = ((~g20876));
assign g24517 = ((~g23822)&(~g22701));
assign II29629 = ((~g21060));
assign g16413 = (g5954&g12075);
assign g8090 = ((~g2944));
assign g27116 = ((~II35301));
assign g13431 = ((~II20592));
assign II37824 = ((~g28386))|((~II37822));
assign g12772 = ((~II19836));
assign II37095 = ((~g28124));
assign II25114 = ((~g18983));
assign g19585 = (g692&g18757);
assign II24299 = ((~g6209))|((~II24298));
assign g7763 = ((~g2394));
assign gbuf156 = (g1954);
assign g10535 = (g7303&g2670);
assign II24156 = ((~g14322))|((~g9407));
assign g27773 = (g5732&g27484);
assign g22610 = (g660&g21473);
assign g16051 = (g12235&g10901);
assign g19781 = (g4535&g17682);
assign g14766 = ((~II21304));
assign II19226 = ((~g10606));
assign g15722 = ((~g13011));
assign g30357 = ((~II39886));
assign II31310 = ((~g22299));
assign g5788 = (g1706&g1760);
assign g22386 = ((~g20837));
assign g6293 = ((~g976));
assign g11249 = ((~II18175));
assign g5711 = (g325&g394);
assign g29810 = (g29748&g22248);
assign g28871 = ((~II37842));
assign g28010 = ((~II36507));
assign II32624 = ((~g17927))|((~g23969));
assign g5748 = (g2400&g2424);
assign g14244 = ((~g12026));
assign g5805 = ((~g243));
assign II16838 = ((~g6945));
assign g5216 = ((~g2667));
assign g7352 = ((~g1148));
assign II40104 = ((~g30342));
assign g18980 = ((~II25031))|((~II25032));
assign g24884 = (g24060&g18917);
assign II31526 = ((~g23684));
assign g13971 = ((~g8846))|((~g12490))|((~g12478));
assign g30725 = ((~II40465));
assign g8537 = (g3410&g960);
assign g14737 = ((~II21286));
assign II14559 = ((~g1735));
assign g12811 = ((~II19872));
assign g10571 = (g7162&g5167);
assign g9785 = (g5473&g1095);
assign g17084 = (g7629&g13954);
assign II27098 = ((~g19199));
assign g20683 = ((~g20198))|((~g3410));
assign g29477 = (g21580&g29275);
assign g15658 = (g8177&g13264);
assign g20332 = ((~g17360));
assign II22014 = ((~g11730));
assign g18973 = ((~g15771));
assign g18567 = ((~g16058)&(~g14551));
assign g22577 = (g13907&g21429);
assign II23498 = ((~g13512));
assign II25710 = ((~g2124))|((~g18048));
assign II25395 = ((~g18782));
assign II27023 = ((~g19550));
assign g16427 = (g5970&g12104);
assign II33000 = ((~g24949));
assign g26706 = ((~II34725));
assign g6022 = ((~g1585));
assign g13151 = ((~g9184));
assign II30847 = ((~g22103));
assign g4985 = ((~g2384));
assign g17585 = ((~II23673));
assign II14786 = ((~g1520));
assign II25781 = ((~g1444))|((~g18207));
assign g8532 = (g6314&g207);
assign g24587 = ((~II32153));
assign g8403 = ((~II15605));
assign g28261 = ((~II37032));
assign II16134 = ((~g6099));
assign g6222 = ((~g2753));
assign g13101 = ((~g9128));
assign II29881 = ((~g21385));
assign g27199 = ((~II35434));
assign II20131 = (g8313&g7542&g2888&g7566);
assign g29499 = ((~II38817));
assign g21005 = ((~g19827)&(~g17875));
assign II32297 = ((~g23968))|((~II32295));
assign g13140 = ((~g9968))|((~g7426));
assign II34343 = ((~g25194));
assign gbuf71 = (g826);
assign g4401 = ((~g1559));
assign g28256 = ((~II37017));
assign II18608 = ((~g10126));
assign g13408 = ((~II20523));
assign g9879 = ((~II16873));
assign g26583 = ((~g25289)&(~g24569));
assign II24326 = ((~g14124))|((~II24325));
assign g20083 = ((~g17968));
assign II29366 = ((~g20966));
assign g28077 = ((~II36676));
assign II31754 = ((~g23712));
assign II35383 = ((~g26160));
assign II25258 = ((~g16974));
assign g7604 = ((~g471));
assign g19420 = ((~II25862));
assign g21804 = ((~g20255))|((~g6838));
assign II15938 = ((~g3338));
assign g28882 = ((~II37851));
assign g20776 = ((~II27365));
assign II18058 = ((~g6643));
assign II33603 = ((~g24519));
assign II36780 = ((~g27577))|((~II36779));
assign II24588 = ((~g9488))|((~II24586));
assign g7192 = ((~g966));
assign g12085 = ((~g11428));
assign g29844 = ((~g29670));
assign g28266 = ((~II37047));
assign II39853 = ((~g30275));
assign g29762 = ((~g16432)&(~g29625));
assign g30941 = ((~II41047));
assign g22587 = (g13927&g21441);
assign II40021 = ((~g30252));
assign II36087 = ((~g27483));
assign g22839 = ((~II29638));
assign g10176 = ((~II17140));
assign g8779 = ((~II15975));
assign g17045 = (g8071&g15474);
assign II26571 = (g18611)|(g18578)|(g18531);
assign II37471 = ((~g27761));
assign g19491 = ((~g17219));
assign II23888 = ((~g14685));
assign g16679 = ((~g14797)&(~g14895));
assign II19563 = ((~g10664));
assign g26381 = (g4951&g25675);
assign g13700 = ((~g13257));
assign II35809 = ((~g26785));
assign g29611 = ((~g13913)&(~g29255));
assign g18966 = ((~g15747));
assign g12256 = ((~II19429));
assign g4421 = ((~g2229));
assign g7895 = ((~II15205))|((~II15206));
assign g19829 = (g18155&g16098);
assign g25375 = (g24683&g18307);
assign g19899 = (g16520&g16895&g16507);
assign g28523 = ((~g26035)&(~g27732));
assign g22213 = ((~g21917));
assign II15505 = ((~g7963));
assign II21458 = ((~g13050));
assign g19598 = (g3925&g17345);
assign g28721 = ((~g28490));
assign g29225 = (g15366&g28785);
assign g19498 = ((~g16767));
assign gbuf217 = (g2700);
assign g14175 = ((~g11980));
assign g16200 = (g5764&g11868);
assign g12173 = ((~g8363));
assign II32368 = ((~g18038))|((~g24012));
assign g13846 = (g7460&g12645);
assign g7626 = ((~g315));
assign g22767 = ((~II29519));
assign g16424 = (g5967&g12101);
assign g30369 = ((~II39916));
assign II30266 = ((~g22744));
assign g13563 = ((~g12711))|((~g3722));
assign g30948 = (g30929&g20786);
assign g22132 = ((~g21395)&(~g19713));
assign g26324 = (g4743&g25579);
assign g19110 = ((~II25303));
assign g5694 = ((~g1681));
assign g13165 = ((~g8305))|((~g3774));
assign II18719 = ((~g8852));
assign g20616 = ((~II27173));
assign g18085 = ((~g16085)&(~g6363));
assign g15556 = (g4939&g12854);
assign II28072 = ((~g19987));
assign g12329 = ((~g10644)&(~g10675)&(~g10692));
assign g19744 = (g17927&g16040);
assign II18142 = ((~g3410));
assign II27711 = (g19262&g19414&g19386);
assign g30543 = ((~II40209));
assign g23882 = ((~II31144));
assign g19836 = (g7143&g18908);
assign g19149 = ((~g17339)&(~g15020));
assign II17963 = ((~g6574));
assign g30755 = (g30632&g22314);
assign g28671 = (g27962&g12161);
assign g28039 = ((~II36574));
assign g26947 = ((~g25798))|((~g26417));
assign g20467 = ((~g17868));
assign gbuf203 = (g2644);
assign II18458 = ((~g11208));
assign II23065 = ((~g9277))|((~g14123));
assign g13286 = ((~g11481)&(~g11332)&(~g11190)&(~g7880));
assign g23632 = (g4171&g22533);
assign g17776 = ((~II23851));
assign II22064 = ((~g12988))|((~II22062));
assign II27984 = ((~g19987));
assign g4144 = ((~g1114));
assign II35678 = ((~g27129));
assign g13819 = ((~g12449));
assign g28327 = (g27900&g22275);
assign II17653 = ((~g6304));
assign g23173 = ((~II29972));
assign g29430 = ((~II38671));
assign II30575 = ((~g23123));
assign II34464 = ((~g25199));
assign g20878 = ((~g19600)&(~g17395));
assign II22973 = ((~g9174))|((~II22972));
assign g28284 = ((~II37101));
assign g8520 = (g6369&g882);
assign II37611 = ((~g28382));
assign II39264 = ((~g29699));
assign II35714 = ((~g26859))|((~g26865));
assign g28940 = (g14207&g28647);
assign g13946 = ((~g12814));
assign g14883 = ((~II21340));
assign II32645 = ((~g18155))|((~g24093));
assign g27503 = ((~II35859));
assign g28735 = ((~g14957)&(~g28430));
assign g23673 = (g17842&g22996);
assign g28060 = ((~II36627));
assign II18007 = ((~g6519));
assign g15528 = ((~II21787));
assign g26853 = (g5716&g26063);
assign II29080 = ((~g21765));
assign g19132 = ((~II25325));
assign g9149 = ((~II16453));
assign g13736 = ((~g13275));
assign g5758 = (g331&g396);
assign g28290 = ((~II37119));
assign II33009 = ((~g24879));
assign II27264 = ((~g19358));
assign II20504 = ((~g11264))|((~g11189));
assign II38820 = ((~g29313))|((~g15933));
assign g24390 = ((~II31844));
assign II21871 = ((~g11718));
assign II26564 = (g18679&g18699&g18728);
assign II38931 = ((~g29209));
assign g23675 = ((~II30823));
assign g25389 = ((~g25005)&(~g5741));
assign g17405 = ((~II23493));
assign g25470 = (g24479&g20400);
assign g24490 = ((~g23686)&(~g22607));
assign g19554 = (g7993&g17240);
assign g10625 = (g7195&g1988);
assign II34316 = ((~g25191));
assign g20279 = ((~g17240));
assign g16240 = (g5804&g11891);
assign g5958 = ((~II14424));
assign g16682 = ((~g14797));
assign II34083 = ((~g25214));
assign g26747 = ((~II34848));
assign g27222 = ((~II35503));
assign g13074 = ((~g9676))|((~g6980));
assign g9764 = (g6448&g411);
assign II13194 = ((~g1315));
assign g18520 = ((~g16171)&(~g14483));
assign II33324 = ((~g25009));
assign II31718 = ((~g23580));
assign g27259 = ((~g26978)&(~g26258));
assign g20382 = ((~g17500));
assign g25291 = ((~g24941));
assign g29484 = (g21544&g29287);
assign g17304 = ((~II23392));
assign g5814 = ((~g927));
assign II16656 = ((~g6066));
assign g12797 = ((~g8350)&(~g8406)&(~g8446));
assign g27515 = ((~II35879));
assign II32633 = ((~g18131))|((~g23970));
assign g24002 = ((~g22812))|((~g14355));
assign g22829 = ((~g21214));
assign II26679 = ((~g17959));
assign g19802 = (g672&g18891);
assign g24823 = ((~II32410))|((~II32411));
assign g15770 = (g5342&g13329);
assign g13953 = (g7646&g12882);
assign II20823 = ((~g13135));
assign II37068 = ((~g28083));
assign g25117 = (g23444&g10974);
assign II23377 = ((~g15763));
assign g24168 = ((~g22400));
assign II30251 = ((~g22628));
assign g17900 = (g4899&g15528);
assign g12883 = ((~g10038)&(~g6284));
assign g13517 = (g5950&g11656);
assign g11710 = ((~g9822))|((~g3678));
assign g28817 = ((~II37778));
assign g24997 = ((~g23528))|((~g1448));
assign II27577 = ((~g20375));
assign g10374 = (g5473&g4775);
assign II26413 = ((~g16643));
assign g11886 = ((~g11126));
assign g29514 = ((~II38872));
assign g10366 = (g6643&g599);
assign g9384 = ((~II16587));
assign g22586 = ((~II29154));
assign g25150 = ((~II32928));
assign g9041 = ((~II16360));
assign II15869 = ((~g7976));
assign g5629 = ((~II14083));
assign g12979 = ((~g9019));
assign II35829 = ((~g26806));
assign g6055 = ((~II14544));
assign g11913 = ((~g11173));
assign g4266 = ((~g1535));
assign II19774 = ((~g10500));
assign II22954 = ((~g14206))|((~II22952));
assign g26311 = (g25911&g9607);
assign II32946 = ((~g24593));
assign g26845 = (g5664&g26056);
assign g28382 = ((~II37291));
assign g23231 = ((~II30146));
assign g27400 = ((~g27012))|((~g6713));
assign g26005 = ((~II33867));
assign g26984 = (g23335&g26558);
assign g11706 = ((~g10928));
assign g10320 = (g7358&g4696);
assign II34159 = ((~g25964));
assign II25579 = ((~g780))|((~II25578));
assign g19981 = (g17729)|(g18419)|(II26429);
assign g18974 = ((~g15774));
assign g8558 = (g7085&g2345);
assign g26050 = ((~g25697)&(~g24922));
assign g9215 = ((~II16489));
assign g29284 = (g29001&g28871);
assign II23866 = ((~g15151));
assign g12293 = ((~g10587)&(~g10628)&(~g10662));
assign g29465 = (g29191&g8424);
assign g12786 = ((~II19847));
assign II18368 = ((~g4325))|((~g4093));
assign g12893 = ((~g8474)&(~g8492)&(~g8508));
assign g29919 = ((~g29736)&(~g22367));
assign g20507 = ((~g18351));
assign g28665 = (g27827&g22222);
assign g29136 = ((~II38151));
assign II31481 = ((~g23556));
assign g21334 = (g9310&g20330);
assign g27407 = (g17914&g27136);
assign II27419 = ((~g19457));
assign g26740 = ((~II34827));
assign g22091 = ((~g21353)&(~g19638));
assign g29631 = ((~II39011));
assign g13176 = ((~g9368));
assign g7925 = ((~g3058));
assign g11870 = ((~g9785)&(~g9910)&(~g10046));
assign g21440 = (g15118&g20424);
assign gbuf60 = (g568);
assign g29557 = (g28789&g29388);
assign g29002 = ((~II37965));
assign g16671 = ((~g14724)&(~g12494));
assign g22157 = ((~g21811))|((~g21816));
assign g29042 = ((~II37999));
assign g15667 = ((~II21918));
assign II24744 = ((~g6167))|((~II24743));
assign g29322 = ((~II38491));
assign g21313 = (g9232&g20311);
assign g19735 = (g17903&g16035);
assign g28274 = ((~II37071));
assign g10471 = (g7265&g2516);
assign g12163 = ((~II19342));
assign II18067 = ((~g6369));
assign g13080 = ((~g9968))|((~g7426));
assign II16228 = ((~g7015));
assign g13108 = ((~g9968))|((~g7426));
assign g28351 = ((~g15605)&(~g28058));
assign g21357 = (g9407&g20356);
assign g24580 = (g18639&g23441&g20043);
assign g5159 = ((~g1272));
assign II37182 = ((~g27791));
assign g27322 = ((~g27070)&(~g26422));
assign g5396 = ((~II13904));
assign II39892 = ((~g30286));
assign g21355 = (g9613&g20354);
assign gbuf64 = (g535);
assign g11523 = ((~II18545));
assign gbuf139 = (g1746);
assign g22603 = ((~II29183));
assign g7996 = ((~g486));
assign g21084 = ((~g20011)&(~g20048));
assign g19290 = ((~II25606))|((~II25607));
assign g13450 = ((~II20649));
assign g8673 = ((~II15869));
assign g26447 = (g5182&g25793);
assign g13446 = ((~II20637));
assign g9524 = ((~II16677));
assign II32661 = ((~g23998))|((~II32659));
assign II30870 = ((~g14194))|((~II30868));
assign g26593 = ((~g25615));
assign g27104 = (g5246&g26466);
assign g27335 = ((~g27087)&(~g26450));
assign g24969 = ((~g23489));
assign g11540 = ((~II18596));
assign g25018 = ((~g23644))|((~g6448));
assign II22025 = ((~g11617));
assign g28460 = (g18091&g27942);
assign g17016 = ((~II22973))|((~II22974));
assign g26427 = (g5118&g25758);
assign g25790 = ((~II33627));
assign g16626 = ((~II22671));
assign g17064 = ((~II23056))|((~II23057));
assign II37323 = ((~g27865))|((~II37322));
assign II28380 = (g20326)|(g18718)|(g18690);
assign g30241 = ((~g30033));
assign g24316 = ((~II31622));
assign II17724 = ((~g6942));
assign g7484 = ((~g2559));
assign II27992 = ((~g20025));
assign g16452 = (g5988&g12156);
assign g10499 = (g5473&g5044);
assign II14143 = ((~g1706));
assign II38348 = ((~g28874));
assign g8340 = (g6369&g909);
assign g8004 = ((~g1174));
assign II18426 = ((~g3722));
assign g30305 = (g2636)|(g2633)|(g30072);
assign g23668 = ((~II30810));
assign g29144 = ((~II38175));
assign g12102 = ((~g11447));
assign g19687 = (g2714&g18833);
assign g30676 = ((~g16419)&(~g30496));
assign II15433 = ((~g2861));
assign II22630 = ((~g13507))|((~g15978));
assign g27031 = (g23340&g26602);
assign g24952 = ((~g23537));
assign II15815 = ((~g3650));
assign g24153 = ((~g22399));
assign g22921 = ((~g16223)&(~g20866)&(~g21293));
assign II16720 = ((~g3774));
assign g12455 = ((~II19637));
assign g28446 = (g18048&g28165);
assign g8489 = (g6519&g939);
assign II40976 = ((~g30799));
assign II16524 = ((~g6000));
assign g19010 = (g13552&g16337);
assign II30188 = ((~g22684));
assign g28579 = ((~II37494));
assign II28649 = ((~g21843));
assign II32491 = ((~g18131))|((~II32490));
assign g26545 = ((~g13790)&(~g25277));
assign II32392 = ((~g17903))|((~II32391));
assign g21732 = ((~g20493)&(~g7329));
assign g30632 = ((~g6119)&(~g30412)&(~g25366));
assign II21595 = ((~g11691));
assign II29348 = ((~g20962));
assign g21569 = (g17825&g18286&g19843&II28103);
assign g10523 = (g7358&g5092);
assign g29792 = (g29491&g10977);
assign II31709 = ((~g23862));
assign g30622 = ((~g6119)&(~g30412)&(~g25393));
assign g9644 = ((~II16747));
assign II40173 = ((~g30497));
assign g27237 = ((~II35548));
assign g23331 = ((~g22999))|((~g22174));
assign II29741 = ((~g21346));
assign g19734 = (g17815&g16034);
assign II40603 = ((~g30614))|((~g30610));
assign g9583 = (g6519&g8218);
assign II39023 = ((~g29508));
assign g28150 = ((~g27387));
assign II13868 = ((~g2180));
assign g10395 = (g7053&g1967);
assign II29984 = ((~g22671));
assign g12023 = ((~g11351));
assign g26085 = (g1448&g25825);
assign g15399 = ((~II21661));
assign g10814 = ((~g5730)&(~g5768)&(~g5816));
assign II28248 = ((~g14309))|((~II28247));
assign g26084 = ((~g25487)&(~g25513));
assign g26366 = (g4916&g25655);
assign II38749 = ((~g29273));
assign g20809 = (g5712&g19113);
assign g22399 = ((~g21230))|((~g14584))|((~g10735));
assign g12437 = ((~II19591));
assign g29622 = (g29250&g11327);
assign g25821 = ((~II33659));
assign g14524 = ((~g12185));
assign II39276 = ((~g29704));
assign g24619 = ((~II32203));
assign g28032 = ((~II36557));
assign II16114 = ((~g7936));
assign II25225 = ((~g16514));
assign II32419 = ((~g24043));
assign g22675 = ((~II29317));
assign g15758 = ((~g12565))|((~g6232));
assign g16293 = ((~g13025));
assign II28435 = ((~g19358));
assign g8525 = (g6783&g1642);
assign g21631 = (g18048&g18474&g19907&II28162);
assign g12980 = ((~g9022));
assign II36096 = ((~g27503));
assign g7830 = ((~g1166));
assign g11441 = ((~II18405));
assign II26472 = (g18635&g18605&g18568);
assign g4076 = ((~g2225));
assign g10726 = ((~g3710))|((~g7358));
assign g12145 = ((~g10364)&(~g10431)&(~g10492));
assign II23920 = ((~g15950));
assign g21849 = (g20272)|(g18651)|(II28374);
assign g26417 = ((~g25969)&(~g24515));
assign II23265 = ((~g9857))|((~II23264));
assign g27263 = ((~g26982)&(~g26269));
assign II39689 = ((~g30035))|((~g30034));
assign II27134 = ((~g19573));
assign II40778 = ((~g30805));
assign II40748 = ((~g30664));
assign g21694 = ((~g20526)&(~g18447));
assign g17093 = ((~II23094))|((~II23095));
assign g12848 = ((~g11059));
assign II23692 = ((~g13540));
assign g6226 = ((~g2818));
assign g30329 = ((~II39828));
assign g14015 = ((~g11897));
assign g29387 = ((~g29019));
assign II25057 = ((~g14186));
assign g9808 = (g6574&g4061);
assign g5676 = (g337&g353);
assign g13241 = ((~g9958));
assign g25939 = ((~g24784));
assign g28289 = ((~II37116));
assign g10450 = (g7162&g4942);
assign g13468 = ((~II20703));
assign g20223 = ((~g18727));
assign g4225 = ((~g701));
assign g29228 = ((~g28996)&(~g28487));
assign II15636 = ((~g3410));
assign g23586 = (g3990&g22473);
assign g22241 = ((~g20655));
assign II25826 = ((~g17168));
assign g26962 = (g6180&g26178);
assign II24112 = ((~g9569))|((~II24110));
assign gbuf123 = (g1564);
assign g15734 = ((~II21982));
assign g12515 = ((~g10773));
assign g5312 = ((~g2655));
assign g13064 = ((~g9822))|((~g7230));
assign II24633 = ((~g7009))|((~II24632));
assign II36728 = ((~g27330));
assign g5687 = (g1018&g1038);
assign g28641 = ((~g27932));
assign g11693 = ((~g9822))|((~g3678));
assign II29004 = ((~g21722));
assign g10231 = ((~II17203));
assign g22193 = ((~g21522)&(~g19857));
assign II21926 = ((~g13126));
assign g21045 = ((~g19886)&(~g18060));
assign g20162 = (g18486&g9757);
assign g11185 = ((~II18103));
assign II22947 = ((~g14015))|((~II22945));
assign g25190 = (g24982)|(g24933);
assign g13385 = (g5815&g11441);
assign g10158 = ((~II17122));
assign II21989 = ((~g11728));
assign g23246 = ((~II30191));
assign g26350 = (g4862&g25620);
assign g9953 = (g7085&g4185);
assign g25984 = ((~II33804));
assign g27443 = ((~II35783));
assign g11786 = ((~II18962));
assign g18948 = ((~g15682));
assign g24428 = ((~g23544)&(~g22398));
assign g15243 = (g7849&g12692);
assign g8068 = ((~g833));
assign g15952 = ((~g11653));
assign g19889 = (g2912&g18943);
assign II21337 = ((~g12408));
assign g26950 = ((~g26417));
assign g23640 = ((~II30776));
assign g10638 = (g7391&g5272);
assign II26651 = (g14936&g18772&g18815);
assign g12077 = ((~g11417));
assign g23819 = ((~II31036))|((~II31037));
assign g26760 = (g26137&g22256);
assign g20120 = ((~g16529)&(~g16924));
assign g20386 = ((~g17517));
assign II34644 = ((~g26159));
assign g29627 = ((~II38999));
assign g17560 = ((~II23648));
assign g15680 = (g5255&g13278);
assign g10448 = (g6980&g4936);
assign II39870 = ((~g30280));
assign g12548 = ((~II19718));
assign g14091 = ((~g11940));
assign g12098 = ((~g10302)&(~g10379)&(~g10444));
assign II35897 = ((~g26817));
assign g25969 = ((~g22917))|((~g24555));
assign g12037 = ((~g11358));
assign g19048 = ((~II25207));
assign g9424 = ((~g5469));
assign II33885 = ((~g25180));
assign II25772 = ((~g762))|((~II25771));
assign g21423 = (g9342&g20414);
assign g19691 = (g16841&g10865);
assign g27003 = (g21996&g26572);
assign II18070 = ((~g5720));
assign g19614 = (g1326&g18787);
assign g17837 = (g4794&g15483);
assign g20910 = ((~g19666)&(~g17527));
assign g11208 = ((~II18130));
assign II18596 = ((~g8870));
assign g18247 = ((~II24247));
assign II23679 = ((~g14966));
assign II30356 = ((~g22902));
assign II16581 = ((~g5438));
assign g20099 = ((~II26535));
assign g17281 = ((~g16081));
assign II40310 = ((~g30503));
assign g19268 = (g14478)|(g16554);
assign g5242 = ((~g1303));
assign g26844 = ((~II34993));
assign g30875 = ((~II40877));
assign g3253 = ((~II13155));
assign g26309 = (g4685&g25554);
assign g21544 = ((~g20025));
assign g25199 = ((~g24558)&(~g20127));
assign g30740 = ((~II40504));
assign g23226 = ((~II30131));
assign g26451 = (g25890)|(g25892);
assign g29503 = ((~II38832))|((~II38833));
assign II29252 = ((~g20924));
assign g13670 = ((~g13234));
assign II32991 = ((~g24599));
assign II23371 = ((~g15761));
assign g20348 = ((~g17402));
assign g9790 = ((~II16838));
assign II21894 = ((~g11720));
assign II25888 = ((~g1457))|((~g18453));
assign g6044 = ((~g2276));
assign g17667 = ((~II23751));
assign g5846 = (g2406&g2441);
assign II21979 = ((~g11727));
assign II16711 = ((~g7015));
assign g24242 = ((~g22309)&(~g21177));
assign g24837 = ((~II32444))|((~II32445));
assign g11642 = ((~g10646));
assign g26735 = ((~II34812));
assign g24905 = (g24084&g18941);
assign g29309 = ((~II38462));
assign II25237 = ((~g16849));
assign g25011 = ((~g23644))|((~g5438));
assign II21900 = ((~g13138));
assign g30059 = ((~g29969)&(~g29811));
assign g12432 = ((~II19582));
assign g23281 = ((~II30296));
assign II30068 = ((~g22647));
assign g11810 = ((~g9605)&(~g9723)&(~g9806));
assign II19877 = ((~g8547));
assign II37269 = ((~g28145));
assign g26633 = ((~g25752));
assign g30747 = ((~II40521));
assign g5937 = ((~g1448));
assign g29296 = ((~g28826));
assign g4916 = ((~g1075));
assign g4954 = ((~g1825));
assign g9909 = (g6519&g4139);
assign g22064 = ((~g21329)&(~g19598));
assign g23240 = ((~II30173));
assign II23309 = ((~g16132));
assign g20412 = ((~g17610));
assign g30790 = ((~g30575)&(~g22387));
assign g20956 = ((~g19936));
assign g7635 = ((~g1693));
assign g13997 = (g7664&g12900);
assign II40507 = ((~g30684));
assign g29104 = ((~II38101));
assign g22979 = ((~II29741));
assign g24368 = ((~II31778));
assign g6102 = ((~II14621));
assign g17352 = (g3942&g14960);
assign g25543 = ((~II33371));
assign II33257 = ((~g24909));
assign g18931 = ((~g15615));
assign II39991 = ((~g30247));
assign g22696 = ((~II29360));
assign g21125 = ((~II27684));
assign II27332 = ((~g19420));
assign II23454 = ((~g15810));
assign II29841 = ((~g21316));
assign II17942 = ((~g5548));
assign II29215 = ((~g20913));
assign g28920 = ((~g28662)&(~g13322));
assign II21629 = ((~g13065));
assign g11231 = ((~II18157));
assign II20583 = ((~g13389));
assign g22245 = (g21690&g12201);
assign g10518 = (g7195&g5081);
assign g15264 = (g1326&g12705);
assign g26611 = ((~g25678));
assign g26506 = ((~II34476));
assign g13237 = ((~g9913));
assign g26647 = ((~g25814));
assign g18812 = ((~g15139));
assign II21694 = ((~g13105));
assign g14797 = ((~g12080));
assign g29610 = (g29349&g11123);
assign g18190 = ((~g14177));
assign g20582 = ((~II27071));
assign II31940 = ((~g24088));
assign II25183 = ((~g18996));
assign g25585 = ((~II33408));
assign g21708 = ((~II28235));
assign g4451 = ((~g2854));
assign g19207 = ((~II25442));
assign g14328 = (g7763&g12997);
assign g5979 = ((~II14449));
assign II30218 = ((~g22794));
assign g26014 = ((~II33894));
assign g30803 = ((~II40661));
assign II36270 = ((~g27549))|((~g15890));
assign g30377 = ((~II39936));
assign gbuf142 = (g1761);
assign II20828 = ((~g13175));
assign II33873 = ((~g25834));
assign g24403 = ((~II31883));
assign II18115 = ((~g8181))|((~II18113));
assign g23555 = ((~II30611));
assign g16044 = ((~g12772));
assign g26654 = ((~g25847));
assign g30629 = ((~g6119)&(~g30412)&(~g25378));
assign g8646 = ((~II15836));
assign g13092 = ((~g10805));
assign II23622 = ((~g15849));
assign II27185 = ((~g20478));
assign g12558 = ((~g8714));
assign g28051 = (g27595&g10021);
assign g17673 = (g4517&g15340);
assign g7562 = ((~g2888));
assign g18024 = ((~II24054))|((~II24055));
assign g24353 = ((~II31733));
assign g16485 = ((~II22557));
assign II39145 = ((~g29613));
assign II15771 = ((~g6000));
assign II32877 = ((~g24567));
assign II35347 = ((~g26265));
assign g24858 = (g24047&g18873);
assign II15466 = ((~g3243));
assign g24521 = ((~g15475)&(~g23859));
assign g18616 = ((~g15074));
assign g8703 = (g6486&g7819);
assign II34121 = ((~g25224));
assign g28125 = ((~II36800));
assign g26349 = ((~II34306));
assign g16012 = ((~g12654));
assign g11643 = ((~g11481)&(~g8045)&(~g7928)&(~g11069));
assign g30502 = (g30199&g11453);
assign g22027 = ((~g21290)&(~g19553));
assign g20221 = (g16825&g10099);
assign g24249 = ((~g22337)&(~g21197));
assign g21432 = ((~g20502)&(~g13335));
assign g4479 = ((~g587));
assign g18636 = ((~g13602));
assign g8651 = ((~II15843));
assign g22332 = ((~g20796));
assign II30751 = ((~g22073));
assign II36987 = ((~g28033));
assign g13162 = ((~g9260));
assign g30090 = (g29840&g11176);
assign II18650 = ((~g8905));
assign g16461 = (g5999&g12176);
assign g5914 = ((~g2185));
assign g21820 = (g16590)|(g19090)|(g16535)|(II28351);
assign g26710 = ((~II34737));
assign g16909 = (g6908&g15033);
assign g25932 = ((~g25125)&(~g17001));
assign gbuf4 = (g2867);
assign g28295 = ((~II37134));
assign g28091 = ((~II36708));
assign II37104 = ((~g28021));
assign g19766 = (g672&g18871);
assign g16100 = (g12130&g10937);
assign g5777 = ((~g1603));
assign g14033 = ((~g12858));
assign II13993 = ((~g2466));
assign g14221 = ((~g12000));
assign II33338 = ((~g25021));
assign g10485 = (g6448&g5024);
assign II14739 = ((~g826));
assign II13947 = ((~g391));
assign g30475 = (g30167&g11315);
assign II30098 = ((~g22711));
assign g8261 = ((~II15451));
assign g28829 = ((~II37790));
assign g21025 = ((~g19860)&(~g17965));
assign g8287 = ((~g3493));
assign II33289 = ((~g25106));
assign II15460 = ((~g3241));
assign g12486 = ((~g8278))|((~g6448));
assign II35893 = ((~g26816));
assign g9605 = (g6574&g8230);
assign II36800 = ((~g27347));
assign g25958 = ((~g22847))|((~g24530));
assign g11923 = ((~II19105));
assign g29393 = ((~g29046));
assign g30931 = ((~g30743)&(~g30750));
assign g28161 = ((~g27428));
assign II18420 = ((~g7015));
assign g20453 = ((~g17785));
assign II25177 = ((~g18985));
assign II24144 = ((~g16278));
assign g24445 = ((~g23427)&(~g22777));
assign g8053 = ((~g141));
assign g8497 = (g3722&g2303);
assign g16794 = ((~II22775));
assign II31074 = ((~g22169));
assign g27185 = (g26126&g22230);
assign g22637 = (g20841&g10927);
assign g25224 = ((~g24772)&(~g23582));
assign g12123 = ((~II19303));
assign g15218 = (g4404&g13180);
assign g10406 = (g7265&g2507);
assign g26302 = (g25903&g9585);
assign g30295 = ((~g13485)&(~g29991));
assign g29939 = ((~g16102)&(~g29792));
assign g20497 = ((~g5410))|((~g18886));
assign g9869 = (g7085&g4076);
assign II25816 = ((~g17162));
assign g30639 = ((~g16186)&(~g30436));
assign g11031 = ((~II17942));
assign g29363 = ((~g28889));
assign g23842 = (g18207&g23041);
assign g24089 = ((~g22922))|((~g14520));
assign g21527 = (g7134&g20468);
assign II33558 = ((~g24460));
assign g23908 = ((~g22353));
assign g20615 = ((~II27170));
assign g5936 = ((~g954));
assign II23415 = ((~g15789));
assign g10765 = ((~g6048));
assign g27564 = ((~g26767)&(~g25184));
assign g27272 = ((~g27000)&(~g26300));
assign g13256 = ((~g10052));
assign g20192 = (g16809&g9228);
assign g29348 = (g1942)|(g1939)|(g29113);
assign g21795 = ((~II28314));
assign g17269 = ((~g16067)&(~g16100));
assign g28874 = ((~g28657)&(~g16221));
assign II18274 = ((~g5837));
assign g23859 = (g22958&g9787);
assign g20754 = ((~II27343));
assign g7228 = ((~g1939));
assign II20529 = ((~g13319));
assign g30717 = ((~II40441));
assign g30317 = ((~II39794));
assign g22686 = (g14124&g21554);
assign g30559 = ((~II40257));
assign II26525 = (g18656&g18670&g18692);
assign II25120 = ((~g18869));
assign II35703 = ((~g26874))|((~II35701));
assign g26627 = ((~g25735));
assign g12000 = ((~g10170)&(~g10257)&(~g10325));
assign g15866 = ((~g12611))|((~g6519));
assign II15226 = ((~g474));
assign II14459 = ((~g805));
assign g11685 = ((~g9822))|((~g3678));
assign g19745 = (g4389&g17601);
assign g26303 = (g25907&g9588);
assign g20182 = (g16705&g16913&g16686);
assign g12692 = ((~II19784));
assign g26773 = (g26145&g22303);
assign g30211 = ((~g30029));
assign g12933 = ((~g8499)&(~g8512)&(~g8527));
assign g23496 = (g5802&g22300);
assign II33542 = ((~g24459));
assign g13048 = ((~g9676))|((~g7162));
assign g8555 = (g7085&g2264);
assign g26818 = ((~g15407)&(~g26335));
assign g19696 = ((~II26123));
assign g7857 = ((~g3055));
assign g28846 = (g27834&g28608);
assign g25927 = ((~g24965))|((~g6448));
assign g16477 = ((~II22533));
assign g8172 = ((~g2975));
assign II19469 = ((~g10664));
assign g8138 = ((~g829));
assign g6512 = ((~g544));
assign g28422 = (g17640&g28150);
assign g25214 = ((~g24754)&(~g23563));
assign II27068 = ((~g19197));
assign g5379 = ((~g3108));
assign II33405 = ((~g25020));
assign II30341 = ((~g22871));
assign II16867 = ((~g3774));
assign g19313 = ((~II25665))|((~II25666));
assign g19798 = ((~II26237));
assign g4865 = ((~g2444));
assign g23001 = ((~g21473));
assign g21060 = ((~g19910)&(~g18152));
assign II25525 = ((~g18803));
assign g17139 = ((~g13957))|((~g13915));
assign II21598 = ((~g13059));
assign g14529 = ((~g11785));
assign g17468 = ((~II23556));
assign g15579 = ((~g12349));
assign g19441 = ((~g17213));
assign II29154 = ((~g20894));
assign g11901 = ((~g11154));
assign g21725 = ((~II28248))|((~II28249));
assign g10559 = (g6713&g5153);
assign g21069 = ((~g20531));
assign g20757 = ((~II27346));
assign g18758 = ((~g14976));
assign g30820 = ((~II40712));
assign g28319 = (g27855&g22246);
assign II14825 = ((~g1231));
assign g19850 = (g4806&g17839);
assign g8087 = ((~II15350));
assign II38169 = ((~g29091));
assign II40907 = ((~g30741));
assign g3649 = ((~g1690));
assign g24226 = ((~g17022)&(~g22282));
assign II16541 = ((~g5438));
assign II34105 = ((~g25221));
assign II21241 = ((~g13378));
assign II30146 = ((~g22712));
assign g12922 = ((~g8961));
assign g24131 = ((~g22484));
assign g8500 = (g6314&g189);
assign g10496 = (g3366&g5035);
assign g15857 = ((~g12565))|((~g6314));
assign g22902 = ((~II29697));
assign g22874 = (g7587&g21708);
assign II38193 = ((~g29099));
assign g27456 = ((~II35796));
assign II28962 = ((~g21721));
assign II21862 = ((~g11717));
assign g16497 = ((~II22593));
assign g21208 = (g20150&g16619&g16586);
assign g10114 = (g6678&g4354);
assign g21269 = (g19681)|(g16797)|(g14936);
assign g22285 = (g21716&g12312);
assign g4708 = ((~g2209));
assign g5186 = ((~g1985));
assign II30206 = ((~g22741));
assign g24377 = ((~II31805));
assign g20725 = ((~II27314));
assign g23267 = ((~II30254));
assign II20745 = ((~g13399))|((~II20743));
assign g30151 = ((~g30014));
assign g27524 = ((~g26931)&(~g24675));
assign g30710 = ((~II40420));
assign II36990 = ((~g28054));
assign g5981 = ((~g207));
assign g22141 = ((~g21401)&(~g19727));
assign II30642 = ((~g22039));
assign g19157 = ((~g17428)&(~g15171));
assign II16085 = ((~g6080));
assign g11906 = ((~g9924)&(~g10060)&(~g10151));
assign g24058 = ((~g22812))|((~g14086));
assign g18225 = ((~II24227))|((~II24228));
assign g10334 = ((~II17300));
assign g20641 = ((~II27232));
assign g6310 = ((~g3101));
assign g9913 = ((~II16915));
assign II29909 = ((~g23050));
assign II20610 = ((~g11812));
assign II40272 = ((~g30366));
assign g23002 = ((~g21477));
assign g22000 = ((~g21268)&(~g19545)&(~g19547));
assign II18791 = ((~g9084));
assign g13182 = ((~g8761)&(~g8778)&(~g8797));
assign II14052 = ((~g870));
assign g28113 = ((~II36766));
assign g29829 = ((~g29665));
assign g15912 = ((~g12611))|((~g6369));
assign g21412 = (g9569&g20404);
assign II24258 = ((~g16463));
assign g23451 = (g18552&g22547);
assign II14596 = ((~g1839));
assign g29245 = ((~II38342));
assign g27903 = ((~II36354));
assign g16987 = (g7555&g15260);
assign g16031 = (g6227&g11747);
assign II25994 = ((~g16860));
assign II32369 = ((~g18038))|((~II32368));
assign g26398 = ((~II34358));
assign g17847 = ((~II23908));
assign g18258 = ((~II24258));
assign g18165 = (g2883&g16287);
assign g7230 = ((~II14937));
assign II19539 = ((~g10549));
assign g22595 = (g13936&g21449);
assign g21891 = (g19302&g11749);
assign g19859 = (g2727&g17871);
assign II38175 = ((~g29092));
assign g21869 = ((~g18319))|((~g19216))|((~g19226));
assign g16391 = (g5939&g12051);
assign g24510 = ((~g15410)&(~g23830));
assign g23773 = ((~II30973));
assign g11492 = ((~II18452));
assign g21149 = ((~g20015)&(~g19981));
assign g13478 = ((~g12611))|((~g3410));
assign g13238 = ((~g9916));
assign II25773 = ((~g18436))|((~II25771));
assign II23433 = ((~g15806));
assign g9125 = (g5473&g7776);
assign g20308 = ((~g17297));
assign g27178 = (g26110&g22213);
assign g28185 = ((~g27356)&(~g26845));
assign II19526 = ((~g10560));
assign g17408 = (g4049&g15049);
assign II33968 = ((~g25372));
assign II20565 = ((~g12432));
assign g30888 = ((~II40916));
assign g4821 = ((~g1739));
assign g16276 = (g1897&g11913);
assign g25035 = ((~g23748))|((~g5512));
assign g11088 = ((~II17998));
assign g19024 = ((~II25135));
assign g26207 = (g2066&g25463);
assign II33692 = ((~g24537));
assign g13097 = ((~g9968))|((~g7488));
assign II27071 = ((~g19218));
assign g26166 = (g686&g25454);
assign g14301 = ((~g12056));
assign g7667 = ((~g3095));
assign II21452 = ((~g13030));
assign g20445 = ((~g17758));
assign II36159 = ((~g27526));
assign II15822 = ((~g3494));
assign g30601 = ((~g30412)&(~g2604));
assign g19202 = (g17919)|(g17998);
assign II31877 = ((~g23766));
assign II14475 = ((~g3225));
assign g18555 = ((~II24633))|((~II24634));
assign g23133 = ((~g17156)&(~g21210));
assign g26053 = (g758&g25306);
assign II40958 = ((~g30742));
assign II36930 = ((~g28071));
assign g10164 = (g3678&g4409);
assign g20589 = ((~II27092));
assign g16229 = (g3772&g11884);
assign II30317 = ((~g22748));
assign g13416 = ((~II20547));
assign g13490 = (g6027&g12220);
assign II37894 = ((~g28584));
assign g27318 = ((~g27060)&(~g26409));
assign g29165 = ((~II38238));
assign g10749 = ((~g6205));
assign II39139 = ((~g29612));
assign II38810 = ((~g29303))|((~g15904));
assign g28338 = (g28029&g19475);
assign g30527 = ((~II40161));
assign g7477 = ((~g1177));
assign g26409 = (g5075&g25732);
assign g15129 = ((~g12094));
assign g23912 = (g14497&g23087);
assign g27299 = ((~g27033)&(~g26371));
assign g19389 = ((~II25810))|((~II25811));
assign g28611 = ((~II37514));
assign g7462 = ((~g2912));
assign II39041 = ((~g29501));
assign g6048 = ((~II14529));
assign g23032 = ((~g21554));
assign g8294 = ((~g3521));
assign g23789 = (g18091&g23024);
assign II24132 = ((~g14107))|((~II24131));
assign II24727 = ((~g14626))|((~II24725));
assign g15521 = ((~II21780));
assign II36135 = ((~g27525));
assign g5035 = ((~g719));
assign II18482 = ((~g8859));
assign g15422 = (g4668&g12794);
assign II34909 = ((~g26265));
assign g11021 = ((~g6030));
assign g15932 = ((~g12711))|((~g7085));
assign g10223 = (g3566&g4535);
assign II38623 = ((~g29293));
assign II38187 = ((~g29086));
assign g19935 = (g2066&g18972);
assign g17794 = (g7423&g16097);
assign g27064 = ((~g26076));
assign II24764 = ((~g6194))|((~II24763));
assign g23013 = ((~g21097)&(~g19254));
assign II22530 = ((~g14774));
assign II29669 = ((~g21073));
assign g11551 = ((~II18629));
assign g28803 = ((~g28493)&(~g28042));
assign g27776 = ((~II36213));
assign g7682 = ((~g1005));
assign g21245 = (g20299&g14837);
assign g15351 = (g4692&g13202);
assign g8363 = ((~II15565));
assign g21914 = ((~II28432));
assign II15499 = ((~g7911));
assign II29220 = ((~g20915));
assign g4842 = ((~g2110));
assign II35968 = ((~g26795));
assign g22277 = ((~g20719));
assign g16085 = ((~g12883))|((~g633));
assign g7388 = ((~g1660));
assign g23218 = ((~II30107));
assign II14715 = ((~g138));
assign g11219 = ((~II18145));
assign g28754 = ((~g28440)&(~g27931));
assign g25602 = ((~II33427));
assign g22592 = ((~II29168));
assign g18896 = ((~g15477));
assign g24256 = (g22003&g11438);
assign g30338 = ((~g14297)&(~g30225));
assign g29940 = ((~II39418));
assign g30904 = ((~II40964));
assign g16851 = ((~g15781)&(~g13000));
assign II39360 = ((~g29766))|((~II39359));
assign g28209 = ((~II36876));
assign II34770 = ((~g26276));
assign g8667 = ((~II15863));
assign g12520 = ((~g8287))|((~g5473));
assign g18916 = ((~g15553));
assign II36870 = ((~g27955));
assign g19650 = (g4076&g17422);
assign g26210 = ((~II34132));
assign g23628 = ((~II30754));
assign g15563 = ((~II21819));
assign g18911 = ((~g15534));
assign g30351 = (g30199&g8408);
assign g7842 = ((~g1165));
assign g29200 = (g15096&g28751);
assign g11761 = ((~g10912));
assign g12527 = ((~g8605));
assign g30569 = ((~g30406));
assign g10763 = ((~g3866))|((~g7426));
assign II15206 = ((~g2972))|((~II15204));
assign II28949 = ((~g21685));
assign II40487 = ((~g30678));
assign II38064 = ((~g28353));
assign II23278 = ((~g9941))|((~II23277));
assign II37065 = ((~g28063));
assign g13551 = ((~g12711))|((~g3722));
assign II22062 = ((~g12999))|((~g12988));
assign g12450 = ((~II19624));
assign g26875 = ((~II35064));
assign g18155 = ((~II24166));
assign g30771 = ((~II40572))|((~II40573));
assign g24080 = ((~g22922))|((~g14573));
assign g13353 = ((~g11481)&(~g8045)&(~g11190)&(~g11069));
assign g17180 = ((~II23243))|((~II23244));
assign g29159 = ((~II38220));
assign II24382 = ((~g13978))|((~II24380));
assign g18955 = ((~g15707));
assign II37808 = ((~g28637));
assign g25136 = ((~II32886));
assign g18537 = ((~II24595))|((~II24596));
assign g10105 = (g5438&g4343);
assign g10082 = (II17042&II17043);
assign g19591 = (g8230&g17330);
assign g21740 = ((~g20198))|((~g6369));
assign g23564 = (g8221&g22434);
assign g15305 = (g4574&g13193);
assign g26521 = ((~g25331));
assign g27817 = ((~II36280));
assign II37771 = ((~g28567));
assign g6130 = ((~II14641));
assign II32985 = ((~g24579));
assign g20967 = ((~g19766)&(~g17735));
assign g9326 = ((~g5906));
assign II29915 = ((~g23055));
assign g20989 = ((~g19802)&(~g17812));
assign g28176 = (g27349&g10940);
assign II39367 = ((~g29767))|((~g15913));
assign g23270 = ((~II30263));
assign g11240 = ((~II18166));
assign II18758 = ((~g8948));
assign g29319 = ((~II38486));
assign II35360 = ((~g26295));
assign II16605 = ((~g7265));
assign g23825 = (g22954&g9644);
assign g29023 = ((~II37982));
assign g4769 = ((~g1048));
assign II36633 = ((~g27304));
assign g13197 = ((~g9531));
assign g15495 = (g4963&g13224);
assign g16266 = ((~g13092));
assign g23353 = ((~g23046))|((~g22204));
assign II14568 = ((~g1071));
assign g13611 = ((~g12926))|((~g3522));
assign g23763 = (g22865&g17688);
assign g30383 = ((~g30306));
assign g20419 = ((~II26846));
assign II26561 = (g14776&g18720&g13657);
assign g23257 = ((~II30224));
assign II31664 = ((~g23516));
assign g8132 = ((~g170));
assign g16924 = ((~g13589));
assign g20708 = ((~II27297));
assign II23530 = ((~g14885));
assign g7357 = ((~II14973));
assign g4093 = ((~g33));
assign g17791 = ((~II23866));
assign II41093 = ((~g30964));
assign g9119 = (g5438&g7754);
assign g13497 = ((~g12657))|((~g3566));
assign II17783 = ((~g7353));
assign II21045 = ((~g12520));
assign g29189 = ((~II38272));
assign g24148 = ((~g22520));
assign g24474 = ((~g23984))|((~g3650));
assign II21551 = ((~g13048));
assign g25168 = ((~II32982));
assign g23275 = ((~II30278));
assign g28790 = ((~g28478)&(~g27991));
assign II14628 = ((~g1846));
assign II15626 = ((~g7265));
assign g23481 = ((~II30525));
assign g13906 = ((~g11822));
assign g28146 = ((~g27631)&(~g17031));
assign g18839 = ((~g15251));
assign g11079 = ((~II17989));
assign g23862 = ((~II31112));
assign g18938 = ((~g15641));
assign g4800 = ((~g1419));
assign g8622 = ((~II15810));
assign g10055 = (g3522&g4254);
assign g26573 = ((~g13839)&(~g25294));
assign g29099 = ((~II38088));
assign g22106 = ((~g21369)&(~g19665));
assign g17570 = ((~II23658));
assign g21154 = (g20193&g12333);
assign g28221 = ((~II36912));
assign g24289 = ((~II31541));
assign g30287 = ((~g16452)&(~g29983));
assign g11856 = ((~g11079));
assign g10587 = (g7230&g5193);
assign g28402 = (g7785&g27839);
assign g7342 = ((~g3024));
assign g4436 = ((~g2486));
assign g4509 = ((~g1030));
assign g11847 = (g2628&g8667);
assign g29350 = ((~II38539));
assign II40808 = ((~g30769));
assign g27709 = ((~II36138));
assign g5623 = ((~g70));
assign II15169 = ((~g2874))|((~II15167));
assign g22402 = ((~g21569));
assign II22593 = ((~g15876));
assign g19630 = (g4029&g17399);
assign II25618 = ((~g18379))|((~II25616));
assign II25358 = ((~g18678));
assign II39809 = ((~g30311));
assign g9928 = (II16930&II16931);
assign g24556 = ((~II32092));
assign g21098 = (g20223&g12204);
assign II18635 = ((~g8904));
assign g11536 = ((~II18584));
assign g10049 = ((~II17009));
assign g16310 = (g5868&g11948);
assign g23458 = (g18602&g22588);
assign II24400 = ((~g13936))|((~II24399));
assign g12067 = ((~g11407));
assign g15470 = (g4763&g12816);
assign g24385 = ((~II31829));
assign g8256 = ((~g30));
assign g23692 = ((~II30860));
assign g27786 = ((~II36227));
assign g10723 = ((~g3554))|((~g6980));
assign g30645 = ((~g16240)&(~g30444));
assign g12366 = ((~II19526));
assign g12860 = ((~II19921));
assign II39392 = ((~g29769))|((~II39391));
assign II31856 = ((~g23635));
assign g25818 = ((~g25077)&(~g21643));
assign II31213 = ((~g22615));
assign g14753 = ((~II21297));
assign II29036 = ((~g21775));
assign II18028 = ((~g7015));
assign g25269 = (g24648&g8700);
assign g26717 = ((~II34758));
assign II23227 = ((~g14090))|((~II23225));
assign g21300 = (g9232&g20288);
assign g23784 = ((~II30994));
assign II37644 = ((~g28341));
assign II13089 = ((~g563));
assign g27949 = (g4406&g27456);
assign II18235 = ((~g6369));
assign g27025 = (g23344&g26594);
assign g19379 = ((~II25782))|((~II25783));
assign g24238 = ((~g17082)&(~g22312));
assign g10652 = (g3618&g5298);
assign II34385 = ((~g25197));
assign II37426 = ((~g27724));
assign g27038 = ((~g26674)&(~g20640));
assign II32520 = ((~g24071))|((~II32518));
assign II18659 = ((~g8938));
assign g30788 = ((~g30602)&(~g22387));
assign g20228 = ((~II26664));
assign g28088 = ((~g26036)&(~g27249));
assign g30220 = (g30040&g8987);
assign g16185 = (g12308&g11017);
assign g19220 = ((~II25463));
assign g30707 = ((~g14131)&(~g30395));
assign g25834 = ((~II33676));
assign II24133 = ((~g9471))|((~II24131));
assign g26615 = ((~g25691));
assign g17877 = (g2998&g15521);
assign g16109 = (g8277&g11803);
assign g26901 = ((~g25627)&(~g26389));
assign II22475 = ((~g2594));
assign g5406 = ((~II13934));
assign g15092 = ((~II21415));
assign II22893 = ((~g15055));
assign g28760 = ((~g15142)&(~g28453));
assign II32679 = ((~g14165))|((~II32677));
assign II34758 = ((~g26221));
assign II27235 = ((~g19420));
assign g7483 = ((~g1834));
assign g10847 = ((~g5800));
assign g5595 = ((~II14049));
assign g8566 = (g6838&g2279);
assign g10842 = ((~II17689));
assign g22726 = (g3036&g21886);
assign II29378 = ((~g20970));
assign g25357 = ((~g24986)&(~g5651));
assign g23509 = ((~g22209));
assign g24230 = ((~g17047)&(~g22291));
assign g19729 = (g4335&g17563);
assign g25159 = ((~II32955));
assign gbuf212 = (g2617);
assign g12006 = ((~g10175)&(~g10262)&(~g10329));
assign II41111 = ((~g30966));
assign II27761 = (g19411&g19382&g19352);
assign g29090 = ((~g28332)&(~g28334));
assign II30501 = ((~g23039));
assign II22694 = ((~g14753));
assign II24982 = ((~g14347));
assign g20318 = ((~g16686)&(~g16913));
assign g22293 = ((~g20743));
assign g8921 = ((~II16209));
assign II36530 = ((~g27276));
assign g30167 = ((~g30018));
assign g14414 = ((~g12978));
assign g19210 = (g18079)|(g18183);
assign g30585 = ((~II40307));
assign g27674 = ((~II36052));
assign g30375 = ((~II39930));
assign II25204 = ((~g16905));
assign g11612 = (g5881&g8378);
assign II29930 = ((~g22176));
assign II18647 = ((~g8851));
assign g6568 = ((~g1339));
assign g21880 = ((~g13854)&(~g19236));
assign g6063 = ((~II14568));
assign II21377 = ((~g11821));
assign g23117 = ((~g17117)&(~g21188));
assign g25087 = ((~g23731));
assign II25567 = ((~g17186));
assign g15858 = ((~g12565))|((~g6232));
assign II31508 = ((~g23613));
assign g30925 = (g30790&g22380);
assign II30669 = ((~g22045));
assign g29215 = ((~g28935)&(~g28471));
assign g12060 = ((~g10251)&(~g10320)&(~g10396));
assign g17194 = ((~g14233))|((~g14132));
assign g5992 = ((~g2156));
assign II23323 = ((~g15664));
assign II22566 = ((~g14883));
assign g20550 = ((~II26985));
assign II18614 = ((~g11002));
assign g17567 = ((~II23655));
assign II18064 = ((~g6519));
assign g19330 = ((~II25717));
assign II16915 = ((~g3494));
assign II23581 = ((~g13528));
assign g13246 = ((~II20295));
assign g8850 = ((~II16092));
assign g29126 = ((~g28373)&(~g27774));
assign g12510 = ((~g8594));
assign g26456 = (g5210&g25811);
assign g21299 = (g9293&g20287);
assign gbuf44 = (g380);
assign II25751 = ((~g2129))|((~II25750));
assign g20559 = ((~II27002));
assign g20603 = ((~II27134));
assign II21508 = ((~g13040));
assign g18486 = ((~g15804));
assign gbuf186 = (g2427);
assign g6431 = ((~g2631));
assign II35915 = ((~g26818));
assign g25744 = ((~II33573));
assign g28655 = ((~g28018));
assign II30368 = ((~g22695));
assign g11512 = ((~II18512));
assign II27958 = ((~g19987));
assign g10340 = (g3866&g7488);
assign II30071 = ((~g22622));
assign II28084 = ((~g20067));
assign g27846 = ((~II36315))|((~II36316));
assign g10456 = (g7195&g4956);
assign II37086 = ((~g28114));
assign II26910 = ((~g17269));
assign II25683 = ((~g17974))|((~II25681));
assign g9438 = (g3254&g8123);
assign g24113 = ((~g22448));
assign g20476 = ((~g17951));
assign g19197 = ((~II25426));
assign g15824 = ((~g12657))|((~g6574));
assign g24279 = ((~II31511));
assign g29789 = ((~g29489)&(~g29242));
assign II23524 = ((~g15833));
assign g26317 = (g25919&g9626);
assign g23794 = ((~II31014));
assign II36615 = ((~g27299));
assign g21888 = ((~g18606))|((~g19298))|((~g19315));
assign g29984 = (g29873&g8351);
assign g10353 = (g7426&g4731);
assign g26190 = ((~II34096));
assign II27868 = ((~g19144));
assign II23879 = ((~g14001))|((~II23878));
assign II17627 = ((~g7575));
assign g30580 = ((~II40294));
assign g25476 = ((~II33304));
assign g13078 = ((~g9822))|((~g7358));
assign g29543 = (g29215&g29380);
assign g5823 = ((~g1612));
assign g19138 = ((~g16781))|((~g16797));
assign g12973 = ((~g9016));
assign g25334 = (g24644&g17984);
assign g20568 = ((~II27029));
assign gbuf36 = (g290);
assign g16473 = ((~II22521));
assign g26754 = (g14657&g26508);
assign g29490 = (g21580&g29301);
assign g16860 = ((~g15828)&(~g13031));
assign g22835 = (g14559&g21678);
assign II24093 = ((~g15096))|((~II24091));
assign II29572 = ((~g21041));
assign g8357 = ((~II15559));
assign g25384 = ((~g24695));
assign g29459 = ((~II38758));
assign g12999 = ((~II20049))|((~II20050));
assign g25254 = ((~g24831)&(~g23687));
assign II23329 = ((~g15760));
assign g5230 = ((~g2810));
assign II28609 = (g21183&g21168&g21148);
assign g22303 = ((~g20763));
assign g4772 = ((~g1060));
assign g22078 = ((~g21342)&(~g19621));
assign II25047 = ((~g14478));
assign g19117 = (g14691&g16644);
assign II37194 = ((~g27800));
assign g17207 = ((~II23287));
assign g15507 = (g5003&g13225);
assign gbuf111 = (g1168);
assign II28219 = ((~g19471))|((~II28217));
assign g11494 = ((~II18458));
assign II24619 = (g14776&g14837&g16142);
assign g27578 = (g24038&g27177);
assign g26623 = ((~g25717));
assign g9755 = ((~g5431));
assign g20144 = (g16679&g16884&g16665);
assign g14580 = ((~g12250));
assign g22233 = ((~g20637));
assign g16090 = ((~g12822));
assign g19169 = ((~II25374));
assign II36957 = ((~g27993));
assign g18828 = ((~g15207));
assign g30962 = ((~g30958));
assign g25957 = (g24782&g11869);
assign g29757 = ((~g16285)&(~g29615));
assign g17617 = (g4409&g15284);
assign g16071 = (g5604&g11777);
assign g20519 = ((~II26966));
assign II24148 = ((~g7079))|((~g14408));
assign II13604 = ((~g125));
assign g5955 = ((~g198));
assign II34002 = ((~g25490));
assign g7146 = ((~g3013));
assign g5850 = ((~II14298));
assign g26049 = ((~g25629)&(~g24908));
assign II31005 = ((~g22149));
assign II29622 = ((~g21055));
assign g25331 = ((~g21230))|((~g14584))|((~g10735))|((~g24603));
assign g4366 = ((~g847));
assign g12272 = ((~g10541)&(~g10600)&(~g10645));
assign g18174 = ((~g14148));
assign g18189 = ((~II24187))|((~II24188));
assign g19620 = (g3984&g17375);
assign g27201 = ((~II35440));
assign g18669 = ((~g13623)&(~g13634));
assign g7989 = ((~g3191));
assign g16112 = (g5684&g11808);
assign g20866 = ((~g19512));
assign II29966 = ((~g22613));
assign g22882 = ((~g21674));
assign II31898 = ((~g23872));
assign g19663 = (g4127&g17451);
assign g30005 = (g29905&g8478);
assign g21033 = ((~g19872)&(~g18011));
assign g30027 = ((~g29565)&(~g29960));
assign g8541 = (g6783&g1651);
assign II29104 = ((~g20881));
assign g20329 = ((~g17348));
assign g12644 = ((~g8780));
assign g15321 = (g4601&g13195);
assign II22869 = ((~g13608));
assign g21655 = ((~II28184));
assign g9527 = ((~g5508));
assign g23832 = ((~II31062));
assign g4818 = ((~g1727));
assign g8689 = ((~II15887));
assign II17100 = ((~g6098));
assign g21487 = (g9941&g20450);
assign g10304 = (g7162&g4659);
assign gbuf56 = (g570);
assign II40628 = ((~g30602))|((~II40627));
assign II22284 = ((~g13348))|((~II22282));
assign II36221 = ((~g27662));
assign g24414 = ((~II31916));
assign g30659 = ((~g16323)&(~g30464));
assign II16034 = ((~g5396));
assign g11583 = ((~II18725));
assign gbuf9 = (g2827);
assign g17200 = ((~II23274));
assign g30501 = ((~II40091));
assign g27714 = ((~II36153));
assign g13524 = ((~g12611))|((~g3410));
assign II26892 = ((~g17246));
assign g18231 = ((~II24235))|((~II24236));
assign II34254 = ((~g25185));
assign g30652 = ((~g16283)&(~g30453));
assign g24282 = ((~II31520));
assign g12266 = ((~g8455));
assign II23794 = ((~g15151));
assign g16069 = (g5346&g11776);
assign II25898 = ((~g2147))|((~II25897));
assign g8621 = (g6486&g6672);
assign II22741 = ((~g14669));
assign II25913 = ((~g1462))|((~g18025));
assign II23959 = ((~g6513))|((~II23958));
assign g21686 = ((~g20164))|((~g6314));
assign II17701 = ((~g6781));
assign g19484 = ((~g16867));
assign g5546 = ((~g3164));
assign g25462 = ((~II33286));
assign g13535 = ((~g12657))|((~g3566));
assign II18497 = ((~g8860));
assign g20975 = ((~g19777)&(~g15421));
assign g23198 = ((~II30047));
assign g27763 = ((~g27534)&(~g27092));
assign g27495 = (g23945&g27146);
assign g27465 = ((~g26846));
assign g18922 = ((~g15574));
assign g19170 = ((~II25377));
assign g5767 = (g1024&g1055);
assign g29912 = ((~g24676)&(~g29716));
assign g19064 = ((~II25253));
assign II24063 = ((~g9326))|((~II24061));
assign g9074 = (g7303&g2639);
assign g9889 = (g6314&g4101);
assign g21187 = ((~g19113));
assign g6281 = ((~g510));
assign g30409 = (g30134&g11025);
assign g10888 = ((~II17753));
assign g16401 = (g5946&g12063);
assign II22855 = ((~g13588));
assign II38905 = ((~g29197));
assign g24509 = ((~g23789)&(~g22674));
assign g5418 = ((~II13968));
assign g27213 = ((~II35476));
assign g24502 = ((~g23743)&(~g22646));
assign g17099 = ((~II23104))|((~II23105));
assign g20896 = ((~g19634)&(~g17462));
assign g17115 = ((~II23114))|((~II23115));
assign g11843 = ((~g9747)&(~g9869)&(~g9952));
assign g15840 = (g8098&g11620);
assign g21845 = ((~g13631)&(~g19161));
assign g22003 = ((~II28557));
assign g11593 = ((~II18755));
assign g25364 = ((~II33198));
assign II32955 = ((~g24584));
assign g13817 = ((~g13336));
assign II22690 = ((~g14703));
assign g17862 = ((~II23923));
assign g20304 = ((~g17288));
assign g12130 = ((~g10788));
assign g5343 = ((~g2796));
assign g30464 = (g30167&g11249);
assign II23436 = ((~g15832));
assign g27630 = ((~g27066))|((~g3774));
assign g13155 = ((~g8688)&(~g8705)&(~g8722));
assign g20899 = ((~g19647)&(~g17474));
assign g5338 = ((~g2658));
assign g15817 = (g8025&g13373);
assign g11525 = ((~II18551));
assign g28932 = ((~II37901));
assign g28692 = ((~II37623));
assign g28394 = ((~g27869)&(~g22344));
assign g23253 = ((~II30212));
assign g26149 = ((~II34041));
assign g27076 = (g5024&g26393);
assign g4314 = ((~g2530));
assign II25463 = ((~g18868));
assign g5750 = ((~g92));
assign g20321 = ((~g17324));
assign g9933 = ((~II16939));
assign g14213 = (g7739&g12973);
assign g9263 = ((~II16517));
assign g26384 = (g4959&g25681);
assign g22738 = (g14292&g21599);
assign g20291 = (g13714&g16302&II26708);
assign II36382 = ((~g27563));
assign g19700 = (g17815&g16024);
assign g24682 = ((~g23688)&(~g24183));
assign g18091 = ((~g14092));
assign g19927 = (g14316&g18463&II26377);
assign g13573 = ((~g12247));
assign g27394 = (g17802&g27134);
assign II16566 = ((~g5556));
assign g25527 = ((~II33355));
assign g29564 = (g28794&g29393);
assign g26310 = (g4688&g25557);
assign g10172 = (g7085&g4433);
assign II16261 = ((~g6448));
assign g19763 = ((~II26198));
assign g6021 = ((~g1579));
assign g30009 = (g29929&g22357);
assign II39032 = ((~g29537));
assign g16288 = (g12308&g11129);
assign II30086 = ((~g22709));
assign II15523 = ((~g3254));
assign g12901 = ((~II19958));
assign g26437 = (g5156&g25773);
assign g27627 = ((~g27012))|((~g3462));
assign II21271 = ((~g11666));
assign g27560 = ((~II35964));
assign g11944 = ((~g11225));
assign II30176 = ((~g22627));
assign g15389 = (g8246&g12772);
assign g24217 = (g22825&g10999);
assign gbuf77 = (g1137);
assign g12991 = ((~g8536)&(~g8549)&(~g8559));
assign g28501 = (g27738)|(g25764);
assign g30681 = ((~g16448)&(~g30330));
assign g30784 = ((~II40618));
assign g22649 = ((~II29265));
assign II24338 = ((~g6632))|((~g14438));
assign g25174 = ((~II33000));
assign g11729 = ((~g9968))|((~g3834));
assign g25328 = (g24644&g17892);
assign g27381 = ((~II35711));
assign g18407 = ((~g15959));
assign g26881 = ((~II35072));
assign g27656 = (g26796&g11004);
assign g3969 = ((~g1531));
assign g29054 = ((~II38011));
assign g19382 = ((~II25791))|((~II25792));
assign II24307 = ((~g13983))|((~II24306));
assign II19844 = ((~g8533));
assign g13854 = (g5349&g12690);
assign g13886 = ((~g12747));
assign g21477 = ((~II28013));
assign II19401 = ((~g10631));
assign II36644 = ((~g27307));
assign g23767 = ((~II30965));
assign g10805 = ((~g5696)&(~g5739)&(~g5786));
assign II39127 = ((~g29608));
assign II30005 = ((~g22757));
assign g10144 = (g3522&g4380);
assign g9287 = ((~g6638));
assign g12336 = ((~II19503));
assign g11775 = ((~g10940));
assign g8821 = ((~II16037));
assign II38854 = ((~g29170));
assign g11964 = ((~g10093)&(~g10182)&(~g10269));
assign g23428 = (g22789&g19607);
assign g29400 = ((~II38591));
assign g8826 = ((~II16050));
assign g5070 = ((~II13742));
assign g5857 = ((~g538));
assign II22551 = ((~g14745));
assign II37026 = ((~g27998));
assign g4851 = ((~g2205));
assign g13494 = ((~g12565))|((~g3254));
assign g17237 = ((~II23323));
assign g27720 = (g27481&g20652);
assign g10869 = ((~II17724));
assign g22644 = ((~g20850))|((~g20904));
assign g24397 = ((~II31865));
assign g27010 = ((~g26063));
assign II25442 = ((~g18866));
assign g29684 = ((~g29562)&(~g29338));
assign g26075 = (g74&g25698);
assign g26251 = ((~II34207));
assign II33900 = ((~g25869));
assign II24062 = ((~g14207))|((~II24061));
assign II18205 = ((~g7975))|((~II18204));
assign g27357 = ((~II35673));
assign g7670 = ((~g317));
assign g22619 = ((~II29203));
assign g27250 = ((~g26955)&(~g26166));
assign II24684 = ((~g16000));
assign g13296 = ((~II20359));
assign g7426 = ((~II14993));
assign II30790 = ((~g22846))|((~g14079));
assign g15592 = (g5021&g12871);
assign g26822 = ((~g15436)&(~g26352));
assign g5741 = ((~g2138));
assign g29580 = ((~g29403)&(~g17031));
assign g21262 = (g20337&g14991);
assign g22852 = ((~II29653));
assign g28706 = ((~II37665));
assign g20579 = ((~II27062));
assign II21661 = ((~g13098));
assign g21371 = (g9264&g20370);
assign g13266 = (g5628&g11088);
assign g19475 = ((~g16725));
assign II29900 = ((~g23125));
assign g23874 = ((~II31136));
assign g8670 = ((~II15866));
assign g15838 = ((~g12711))|((~g6838));
assign g8718 = ((~II15922));
assign g15624 = (g5186&g13261);
assign g29700 = ((~II39154));
assign II31838 = ((~g23585));
assign II36903 = ((~g28045));
assign II35940 = ((~g26823));
assign g28906 = ((~II37875));
assign g12392 = ((~II19552));
assign gbuf216 = (g2697);
assign g13838 = ((~g13361));
assign g20428 = ((~g17676));
assign II14775 = ((~g823));
assign II17819 = ((~g6448));
assign g18492 = ((~II24538))|((~II24539));
assign II32248 = ((~g23919));
assign g9310 = ((~g5811));
assign g19017 = ((~II25114));
assign g17493 = ((~II23581));
assign g9895 = ((~II16897));
assign g11720 = ((~g9968))|((~g3834));
assign g22473 = ((~II29019));
assign g10414 = (g7426&g4876);
assign II23171 = ((~g9471))|((~g13881));
assign II36999 = ((~g28076));
assign g17397 = (g4023&g15040);
assign II13122 = ((~g20));
assign II39873 = ((~g30281));
assign II38466 = ((~g28754));
assign g15585 = ((~II21841));
assign g29299 = ((~II38440));
assign gbuf199 = (g2625);
assign g27584 = ((~g26938)&(~g24736));
assign g4335 = ((~g162));
assign g5061 = ((~g1407));
assign g5923 = ((~II14381));
assign g9091 = (g3306&g7670);
assign g11961 = ((~g11256));
assign II21560 = ((~g11685));
assign g24121 = ((~g22455));
assign g9487 = ((~II16656));
assign g19029 = ((~II25150));
assign g12443 = ((~II19605));
assign g27684 = ((~II36063));
assign II19582 = ((~g8862));
assign g28173 = ((~g27486));
assign g9795 = ((~g6019));
assign g15030 = (g4110&g13158);
assign g27581 = ((~g26925)&(~g24728));
assign g23745 = ((~II30941));
assign II36539 = ((~g27279));
assign II20832 = ((~g12507));
assign g25185 = ((~g24492)&(~g10024));
assign g7566 = ((~g2896));
assign II17957 = ((~g6713));
assign g24543 = ((~g23891)&(~g22764));
assign g13131 = ((~g9968))|((~g7426));
assign II21825 = ((~g13127));
assign g8562 = (g6783&g1588);
assign g23666 = (g22851&g20407);
assign g29265 = ((~II38379))|((~II38380));
assign g19904 = (g2059&g18949);
assign II26461 = (g18096)|(g17998)|(g17919);
assign g27914 = (g13927&g27404);
assign g16137 = (g12275&g10983);
assign g26023 = (g25422&g24912);
assign II33683 = ((~g24472));
assign g16594 = ((~g15933)&(~g15913)&(~g14650));
assign g8449 = ((~II15651));
assign g17591 = ((~II23679));
assign II24751 = ((~g7455))|((~g14609));
assign g20840 = (g5885&g19132);
assign g23263 = ((~II30242));
assign II13092 = ((~g1249));
assign II28247 = ((~g14309))|((~g19494));
assign g17111 = ((~g14753)&(~g14737)&(~g15952));
assign II38539 = ((~g29113));
assign II27621 = ((~g20417));
assign g13275 = ((~II20334));
assign II25015 = ((~g14158));
assign II16744 = ((~g3338));
assign g25283 = ((~g24929));
assign II14951 = ((~g2619));
assign g11671 = ((~II18857));
assign II31700 = ((~g23835));
assign II33168 = ((~g25042));
assign II24602 = ((~g6890))|((~II24601));
assign g19887 = (g18155&g16179);
assign g18935 = ((~g15631));
assign II40588 = ((~g30629))|((~II40587));
assign g29725 = ((~g29583)&(~g1911));
assign g18128 = (g5187&g15682);
assign g25310 = (g24704&g8813);
assign g28741 = ((~II37702));
assign II17673 = ((~g8107));
assign g10263 = ((~II17225));
assign g5703 = ((~g109));
assign g29656 = ((~II39086));
assign g15737 = ((~g12412));
assign g16056 = ((~g12791));
assign g24863 = ((~g24258))|((~g23319));
assign g20993 = ((~g19807)&(~g17835));
assign II16556 = ((~g7015));
assign II19360 = ((~g10683));
assign II22726 = ((~g14642));
assign g18419 = ((~II24437))|((~II24438));
assign g4006 = ((~g160));
assign II16486 = ((~g5473));
assign g12109 = ((~II19289));
assign g5642 = ((~g61));
assign g17216 = ((~g4495)&(~g14529));
assign g26371 = (g4919&g25658);
assign g11835 = ((~g11039));
assign g13608 = ((~II20828));
assign g19183 = ((~II25402));
assign II18801 = ((~g11331))|((~II18799));
assign g30688 = ((~g13484)&(~g30348));
assign g9098 = (g5512&g7691);
assign g11628 = ((~II18810));
assign II21569 = ((~g11686));
assign II36447 = ((~g27257));
assign g18060 = (g5129&g15647);
assign II16870 = ((~g7265));
assign g17503 = ((~II23591));
assign g10252 = ((~g7802))|((~g3678));
assign g27164 = ((~g26466));
assign II34812 = ((~g26280));
assign II14848 = ((~g2824));
assign II21855 = ((~g13113));
assign g28169 = ((~g27467));
assign g4430 = ((~g2250));
assign g8783 = (g7303&g7865);
assign g22747 = ((~II29475));
assign g27085 = (g22134&g26642);
assign g18474 = ((~g14502));
assign g6313 = ((~II14731));
assign g24539 = ((~II32067));
assign g8711 = ((~II15915));
assign g27276 = ((~g27004)&(~g26316));
assign g21811 = (g19138)|(g16974)|(g14936);
assign II16059 = ((~g3878));
assign II41035 = ((~g30796));
assign g22706 = ((~II29378));
assign g22663 = ((~II29291));
assign II26028 = ((~g16566));
assign g19307 = (g17063&g8587);
assign g26174 = ((~II34074));
assign g19184 = ((~g17798)&(~g15520));
assign g28702 = ((~II37653));
assign g10988 = ((~II17889));
assign g26588 = ((~g25602));
assign g24084 = ((~g23077));
assign II29055 = ((~g21732));
assign g8762 = (g3806&g7892);
assign II15191 = ((~g2956))|((~II15190));
assign g9183 = ((~II16469));
assign g7224 = ((~g1845));
assign II39348 = ((~g29732))|((~II39347));
assign g23357 = ((~g22210)&(~g20127));
assign g11407 = ((~II18365));
assign g23799 = ((~II31021));
assign II25904 = ((~g17194));
assign g28486 = (g18379&g27994);
assign g9870 = (g6838&g4079);
assign g12765 = ((~II19829));
assign II20324 = ((~g10124));
assign g18007 = ((~g14464)&(~g16036));
assign g10297 = (g5473&g4647);
assign g17189 = ((~II23253));
assign II31043 = ((~g22161));
assign II21658 = ((~g13072));
assign g24105 = ((~g22425));
assign g28745 = ((~g28431)&(~g27922));
assign g15853 = ((~g13310))|((~g12354));
assign g29530 = ((~II38898));
assign g24035 = ((~II31257));
assign g4609 = ((~g590));
assign II16958 = ((~g7391));
assign g23041 = ((~g21573));
assign g5976 = ((~II14442));
assign g17162 = ((~g14027))|((~g13971));
assign g21906 = (g5715&g20513);
assign g19667 = (g1319&g18826);
assign II35458 = ((~g26886));
assign g17948 = (g4967&g15566);
assign g21824 = ((~II28357));
assign gbuf18 = (g2854);
assign g20938 = ((~g19721)&(~g17631));
assign g10307 = (g6980&g4668);
assign g20947 = ((~g19734)&(~g15335));
assign g20177 = (g13677&g13750&II26615);
assign g29690 = ((~II39124));
assign g19350 = ((~g17094));
assign g24260 = ((~II31454));
assign g21374 = (g9407&g20373);
assign g8602 = ((~II15794));
assign g24295 = ((~II31559));
assign II27365 = ((~g19401));
assign g12053 = ((~g11382));
assign g24547 = ((~g15639)&(~g23914));
assign g4205 = ((~g131));
assign II22988 = ((~g15296))|((~g14321));
assign g20563 = ((~II27014));
assign g27972 = ((~II36441));
assign g24399 = ((~II31871));
assign g21950 = ((~II28476));
assign g25243 = ((~g24803)&(~g23631));
assign g5201 = ((~g2451));
assign g12436 = ((~g8587)&(~g10749));
assign II19823 = ((~g10705));
assign g19675 = (g2013&g18831);
assign g4558 = ((~g2206));
assign II25171 = ((~g16528));
assign II25790 = ((~g2133))|((~g17954));
assign g18121 = ((~g14402));
assign g26969 = (g23320&g26543);
assign II39647 = ((~g30058));
assign g22009 = ((~g19283))|((~g21179))|((~g19333));
assign g13620 = ((~II20844));
assign g20593 = ((~II27104));
assign g27091 = (g5142&g26429);
assign g27831 = ((~II36296));
assign g13457 = ((~II20670));
assign II21923 = ((~g11722));
assign II20022 = (g9488&g9407&g9342&g9277);
assign II40233 = ((~g30363));
assign g9120 = (g3618&g7757);
assign g24597 = ((~II32175));
assign g30851 = ((~II40805));
assign g19679 = (g4188&g17482);
assign g24333 = ((~II31673));
assign g24220 = ((~g22750));
assign g23325 = ((~g23080))|((~g23070));
assign II40676 = ((~g30640));
assign g26595 = ((~g25623));
assign g25951 = (g24800&g13670);
assign g24054 = ((~g22852))|((~g14374));
assign g25142 = ((~II32904));
assign II40459 = ((~g30669));
assign g25182 = (g24681&g20676);
assign g30865 = ((~II40847));
assign g29450 = ((~II38731));
assign g17992 = ((~II24029))|((~II24030));
assign II32659 = ((~g18038))|((~g23998));
assign g19815 = (g2033&g17770);
assign II33427 = ((~g25044));
assign g20351 = ((~g17413));
assign g14746 = ((~II21292));
assign g22548 = ((~II29098));
assign g11852 = ((~g11063));
assign g4783 = ((~g1265));
assign g23020 = ((~g21524));
assign g23208 = ((~II30077));
assign II32452 = ((~g18038))|((~II32451));
assign g19532 = (g16943)|(g16770)|(g16712);
assign II32615 = ((~g18247))|((~g24091));
assign g16132 = ((~II22283))|((~II22284));
assign II31775 = ((~g23837));
assign g11996 = ((~g11306));
assign g12106 = ((~g11459));
assign g17425 = ((~II23513));
assign g25979 = ((~g24611)&(~g23538));
assign g22032 = ((~g21300)&(~g19559));
assign g3239 = ((~II13113));
assign g17454 = ((~II23542));
assign II33894 = ((~g25868));
assign II18626 = ((~g8649));
assign g19246 = (g18395)|(g18478);
assign g30938 = ((~II41038));
assign II34306 = ((~g25259));
assign g21338 = (g9391&g20335);
assign g23372 = ((~g22000))|((~g21988));
assign g17062 = (g7613&g15544);
assign II30994 = ((~g22147));
assign g18276 = ((~II24272))|((~II24273));
assign II29023 = ((~g20672));
assign g16221 = (g5614&g13257);
assign II38405 = ((~g28723));
assign II37313 = ((~g27883))|((~II37311));
assign g4575 = ((~g2503));
assign II40221 = ((~g30349));
assign g28159 = ((~g27419));
assign II36776 = ((~g27342));
assign g25431 = ((~g24969));
assign g9649 = ((~g5982));
assign g20135 = (g18486&g9885);
assign g18328 = ((~g14768));
assign g21121 = (g20054&g14244);
assign g4512 = ((~g1056));
assign II28956 = ((~g21714));
assign g8175 = ((~II15398));
assign g29380 = ((~g28979));
assign g19059 = ((~II25240));
assign II33411 = ((~g24491));
assign g22557 = (g21907&g12654);
assign II29426 = ((~g20989));
assign g24871 = ((~g16422)&(~g24256));
assign g5908 = ((~g1624));
assign gbuf110 = (g1161);
assign g28049 = ((~II36604));
assign g8510 = (g6574&g1639);
assign g25784 = ((~II33621));
assign g5612 = ((~II14066));
assign g29065 = ((~II38024));
assign g4922 = ((~g1266));
assign g27760 = ((~g27509)&(~g27076));
assign g12187 = ((~g8285));
assign g11730 = ((~g9822))|((~g3678));
assign g29653 = ((~II39077));
assign g27662 = ((~II36042));
assign g27157 = ((~g23471)&(~g26067));
assign II39418 = ((~g29668));
assign g24945 = ((~g23533));
assign g7520 = ((~g2830));
assign g26802 = ((~g26188)&(~g25466));
assign g27043 = (g23349&g26609);
assign II25510 = ((~g18542));
assign II34140 = ((~g25230));
assign g19095 = (g14922&g18765&g16266&g16313);
assign g10464 = (g7358&g4976);
assign g19431 = ((~II25872));
assign g18569 = ((~II24662));
assign g28774 = ((~g28457)&(~g27951));
assign II41064 = ((~g30927))|((~g30926));
assign g24439 = (g14703&g15962&g24153);
assign g8901 = ((~II16179));
assign g10895 = ((~II17768));
assign g16197 = (g518&g11862);
assign II15843 = ((~g3650));
assign g21947 = ((~II28467));
assign g11708 = ((~g9534))|((~g3366));
assign g11955 = ((~g10074)&(~g10165)&(~g10249));
assign g24974 = (g7600&g24030);
assign g26009 = ((~II33879));
assign II34535 = ((~g25451));
assign g4882 = ((~g391));
assign II18557 = ((~g8810));
assign g22900 = ((~g16223)&(~g20956));
assign g20284 = (g18744&g18815&g13774&g16433);
assign g23312 = ((~II30389));
assign II36772 = ((~g27341));
assign g21404 = ((~II27949));
assign g22152 = ((~g21422)&(~g19748));
assign g19237 = ((~II25486));
assign II25132 = ((~g16862));
assign II34473 = ((~g25288));
assign g17500 = ((~II23588));
assign g17485 = (g4089&g16013);
assign g11972 = ((~g11277));
assign g30227 = (g30048&g9058);
assign g12539 = ((~g10408)&(~g10472)&(~g10531));
assign g30301 = ((~g13504)&(~g30002));
assign II20444 = ((~g10869));
assign II24353 = ((~g9356))|((~II24351));
assign g19603 = (g692&g18786);
assign g7263 = ((~g1662));
assign II16590 = ((~g5473));
assign g29562 = (g29228&g29392);
assign II19624 = ((~g9354));
assign g30494 = ((~II40078));
assign II31082 = ((~g22170));
assign II24702 = ((~g7259))|((~g14554));
assign g15257 = (g4357&g12702);
assign II34044 = ((~g25566));
assign g10124 = ((~g5326));
assign g12044 = ((~g10212)&(~g10299)&(~g10375));
assign g26038 = (g25589&g19504);
assign g8965 = ((~II16273));
assign II26154 = ((~g16851));
assign g20052 = (g16804&g3134);
assign g25860 = ((~g24630));
assign g20536 = ((~g18539));
assign g17914 = ((~g13963));
assign g23467 = (g18634&g22625);
assign g12379 = ((~II19539));
assign g16602 = ((~g14565));
assign II21012 = ((~g12503));
assign g6901 = ((~g3006));
assign II16517 = ((~g6000));
assign II19587 = ((~g9173));
assign g27309 = ((~g27049)&(~g26388));
assign II23317 = ((~g16181));
assign g18787 = ((~g15049));
assign g5794 = ((~g2288));
assign g24387 = ((~II31835));
assign g9290 = ((~II16532));
assign II40820 = ((~g30745));
assign g29176 = (g29097&g20690);
assign g29642 = ((~II39044));
assign g24306 = ((~II31592));
assign g23601 = ((~II30701));
assign g8699 = ((~II15899));
assign g29354 = ((~g29127)&(~g17031));
assign II14802 = ((~g551));
assign g13227 = ((~g9880));
assign g28122 = (g27617&g10334);
assign g23626 = ((~II30748));
assign g26231 = (g2760&g25472);
assign II35946 = ((~g14904))|((~II35944));
assign g28026 = ((~II36545));
assign g8023 = ((~II15317));
assign g17782 = ((~II23857));
assign g8486 = (g6314&g261);
assign g9022 = ((~II16344));
assign g26332 = (g4769&g25590);
assign g17510 = (g4231&g15185);
assign g11500 = ((~II18476));
assign g19936 = ((~g16650))|((~g10082));
assign g30829 = ((~II40739));
assign g8861 = (g6643&g493);
assign II15830 = ((~g8031));
assign g24762 = (g12876&g24114);
assign g27208 = ((~II35461));
assign g15870 = ((~g12657))|((~g6783));
assign g24073 = ((~g23059));
assign g19502 = ((~g16775));
assign II15313 = ((~g2930));
assign g15599 = ((~II21855));
assign g28090 = ((~II36705));
assign g15710 = (g5227&g12935);
assign g21105 = ((~g20052)&(~g20088)&(~g20109));
assign g23955 = ((~II31213));
assign g4714 = ((~g2240));
assign II31568 = ((~g24033));
assign g21439 = (g9569&g20423);
assign g27858 = ((~II36327));
assign g24937 = ((~II32687))|((~II32688));
assign g4677 = ((~g1516));
assign g9273 = ((~II16521));
assign g30547 = ((~II40221));
assign II16681 = ((~g6643));
assign g29964 = (g29757&g13786);
assign g12698 = ((~g11347)&(~g11420)&(~g8327));
assign II16598 = ((~g3618));
assign g23294 = ((~II30335));
assign II20100 = (g10186&g3018&g3028);
assign II19377 = ((~g10560));
assign g18583 = ((~g13741));
assign g30348 = (g30203&g8400);
assign g11531 = ((~II18569));
assign g12180 = ((~g10407)&(~g10471)&(~g10530));
assign II32604 = ((~g23339));
assign II32973 = ((~g24572));
assign g27538 = ((~g24982)&(~g24672)&(~g26784));
assign g4752 = ((~g593));
assign II20805 = ((~g13124));
assign g27247 = (g27011&g16702);
assign g20218 = (g16325&g13805&g13825&II26651);
assign g30765 = ((~g30685));
assign g29184 = ((~g28852)&(~g28411));
assign g11572 = ((~II18692));
assign II34677 = ((~g26232));
assign g20952 = ((~g19744)&(~g15349));
assign II15580 = ((~g5837));
assign II15975 = ((~g5744));
assign g27728 = (g27564&g20766);
assign g24379 = ((~II31811));
assign II32356 = ((~g18014))|((~II32355));
assign g26934 = ((~II35124))|((~II35125));
assign II28068 = (g17802&g18265&g17882);
assign II36473 = ((~g27262));
assign g29539 = (g27754&g29377);
assign g13051 = ((~g9822))|((~g7358));
assign g28435 = (g17937&g28160);
assign II38053 = ((~g28350));
assign g27326 = ((~g27074)&(~g26427));
assign g27489 = ((~II35837));
assign g8107 = ((~II15372));
assign g9777 = (g6519&g4032);
assign g5988 = ((~g1570));
assign g13304 = ((~g10266));
assign g23870 = ((~II31124));
assign gbuf53 = (g513);
assign g28270 = ((~II37059));
assign g16217 = (g5776&g11876);
assign II34964 = ((~g26547));
assign g20270 = (g14797&g18692&g13657&g16243);
assign g12113 = ((~g10322)&(~g10399)&(~g10463));
assign g21116 = ((~g20086)&(~g20107)&(~g20131));
assign g23400 = ((~g17540)&(~g22597));
assign g5667 = ((~g222));
assign g24566 = ((~g23944)&(~g22842));
assign II39767 = ((~g30061));
assign g28528 = ((~g26030)&(~g27728));
assign g21955 = ((~II28491));
assign g24320 = ((~II31634));
assign g12816 = ((~II19877));
assign g23571 = (g3931&g22445);
assign g18390 = ((~g14414));
assign g29152 = ((~II38199));
assign g17607 = ((~II23695));
assign g25161 = ((~II32961));
assign g27963 = (g4545&g27467);
assign g9000 = ((~II16318));
assign II40718 = ((~g30654));
assign g7613 = ((~g1158));
assign g19323 = ((~g17059));
assign II24544 = ((~g14263))|((~g9649));
assign g27304 = ((~g27044)&(~g26381));
assign g26977 = (g23320&g26550);
assign II21351 = ((~g12420));
assign II34168 = ((~g25237));
assign g5018 = ((~g2804));
assign II40291 = ((~g30468));
assign g18101 = ((~g14099));
assign g27267 = ((~g26995)&(~g26290));
assign II15961 = ((~g6051));
assign g21017 = ((~g19848)&(~g17926));
assign g28473 = ((~g27730)&(~g26794));
assign g23048 = ((~g21586));
assign g21858 = ((~g18096))|((~g19194))|((~g19202));
assign II37596 = ((~g28377));
assign g25040 = ((~g23923))|((~g6486));
assign g4684 = ((~II13578));
assign g21136 = (g19271&g19261&II27695);
assign g25201 = ((~g24575)&(~g18407));
assign g9904 = (g3366&g4124);
assign II34740 = ((~g26465));
assign g16845 = ((~g15755)&(~g12990));
assign II16021 = ((~g6060));
assign II23570 = ((~g15871));
assign g4386 = ((~g1394));
assign g5292 = ((~g2857));
assign g6115 = ((~II14628));
assign g7577 = ((~g805));
assign g23407 = ((~g17630)&(~g22634));
assign II25506 = ((~g18781));
assign g20572 = ((~II27041));
assign II31266 = ((~g22242));
assign g17321 = ((~II23409));
assign g26650 = ((~g25830));
assign II25881 = ((~g776))|((~II25880));
assign g28660 = (g27916&g11911);
assign II33617 = ((~g24522));
assign g12875 = ((~g10779));
assign g21973 = ((~g21251)&(~g19520));
assign g28407 = (g7799&g27858);
assign g18690 = (g14936&g15080&g13774&g16371);
assign g11017 = ((~II17928));
assign g18908 = ((~g15521));
assign II29307 = ((~g20946));
assign g11930 = ((~g11202));
assign II25761 = ((~g79))|((~g17882));
assign II17922 = ((~g8031));
assign II18124 = ((~g6314));
assign II32687 = ((~g18155))|((~II32686));
assign g26861 = ((~II35028));
assign II39577 = ((~g29939));
assign g13030 = ((~g9676))|((~g7162));
assign g17691 = ((~II23775));
assign g27077 = (g22083&g26636);
assign g4736 = ((~II13604));
assign g20090 = (g18063&g3120);
assign g18804 = ((~g13905)&(~g12331));
assign g16009 = (g12071&g10843);
assign II32310 = ((~g23973))|((~II32308));
assign g9634 = (g6314&g3934);
assign g27280 = ((~g27008)&(~g26325));
assign g16469 = ((~II22509));
assign II28181 = (g14124&g14559&g14222);
assign g20064 = ((~g17209))|((~g2160));
assign g30832 = ((~II40748));
assign II23895 = ((~g9174))|((~II23893));
assign II37410 = ((~g27722));
assign II17904 = ((~g6713));
assign g30393 = (g30233&g8984);
assign g21666 = (g3398&g20504);
assign II19608 = ((~g10831));
assign g21073 = ((~g19928)&(~g18244));
assign g27931 = (g4221&g27432);
assign g19810 = (g17927&g16090);
assign g29735 = ((~g23797)&(~g29583));
assign g8460 = ((~II15662));
assign g10259 = (g3722&g4570);
assign II20646 = ((~g13323));
assign g30973 = ((~II41093));
assign II37071 = ((~g28064));
assign g25021 = ((~g23694))|((~g5473));
assign g20344 = ((~g17384));
assign g13786 = ((~g13300));
assign II33915 = ((~g25762));
assign g19570 = (g8150&g17291);
assign II39939 = ((~g30300));
assign II29320 = ((~g20950));
assign g6033 = ((~g1582));
assign g12214 = ((~g10457)&(~g10518)&(~g10580));
assign g17632 = (g4441&g15311);
assign g29828 = (g29740&g20802);
assign II13179 = ((~g853));
assign g5872 = (g1718&g1764);
assign II19452 = ((~g10560));
assign g25309 = (g5697&g24864);
assign g29865 = ((~g29678));
assign g24965 = (g23922)|(g23945);
assign g28910 = (g28612&g9303);
assign g24783 = ((~g16161)&(~g24224));
assign II30212 = ((~g22742));
assign g5969 = ((~g1642));
assign II35872 = ((~g26925));
assign gbuf143 = (g1763);
assign II24512 = ((~g13992))|((~g9342));
assign g30033 = ((~g24723)&(~g29931));
assign g26666 = ((~g25216)&(~g10133));
assign g20984 = ((~II27531));
assign g27072 = (g22021&g26633);
assign g5773 = ((~g1227));
assign II39384 = ((~g29718))|((~g29710));
assign g13645 = (g6281&g12504);
assign g4110 = ((~g414));
assign g8129 = ((~g151));
assign g11898 = ((~g11145));
assign g26501 = ((~II34469));
assign g30794 = ((~II40640));
assign g15204 = ((~II21494));
assign II32539 = ((~g18247))|((~II32538));
assign g21326 = (g9613&g20325);
assign g26709 = ((~II34734));
assign g15769 = (g5341&g13328);
assign g8509 = (g6783&g1633);
assign g29927 = ((~II39376))|((~II39377));
assign g20461 = ((~g17839));
assign g10927 = ((~g6153));
assign II38940 = ((~g29213));
assign g28193 = (g27573&g21914);
assign g15173 = (g4347&g13177);
assign g13128 = ((~g9822))|((~g7358));
assign II23676 = ((~g15868));
assign g22184 = ((~g21489)&(~g19823));
assign II38947 = ((~g29218));
assign g13009 = (g3995&g10416);
assign g22312 = (g21752&g12349);
assign g29193 = ((~II38282));
assign g16655 = ((~g15933)&(~g14669)&(~g15890));
assign II39249 = ((~g29693));
assign g26048 = ((~g25628)&(~g24906));
assign g30485 = ((~g14098)&(~g30220));
assign g20490 = ((~g18166));
assign g17707 = ((~II23791));
assign g23056 = ((~g21594));
assign g28714 = (g28394&g22306);
assign II28728 = ((~g13519))|((~II28726));
assign g7553 = ((~g3114));
assign g24496 = ((~g23724)&(~g22633));
assign II16182 = ((~g5407));
assign g16027 = ((~g12744));
assign g22089 = ((~g21351)&(~g19632));
assign g7554 = ((~g117));
assign g25049 = ((~g23984))|((~g7195));
assign g9134 = ((~II16438));
assign II31544 = ((~g23438));
assign g7834 = ((~g2953));
assign II24251 = ((~g7329))|((~g14520));
assign g22039 = ((~g21306)&(~g19566));
assign II36454 = ((~g27588));
assign g25195 = (g24993)|(g24945);
assign g26727 = ((~II34788));
assign II24265 = ((~g9232))|((~II24263));
assign g13293 = ((~g10214));
assign g21419 = (g9795&g20409);
assign g10991 = ((~II17892));
assign g11819 = ((~g11014));
assign g25493 = ((~II33321));
assign g11828 = ((~g9639)&(~g9764)&(~g9892));
assign II17916 = ((~g7560));
assign g30817 = ((~II40703));
assign g25562 = ((~II33390));
assign g19910 = (g2746&g18953);
assign g17577 = (g4351&g15251);
assign g28042 = (g14559&g27543);
assign g20111 = (g18261&g9884);
assign II16231 = ((~g5414));
assign II20479 = ((~g10849));
assign II23689 = ((~g15920));
assign II29229 = ((~g20805));
assign g13002 = ((~g8556)&(~g8565)&(~g8572));
assign II35542 = ((~g26858));
assign g13112 = ((~g9534))|((~g6678));
assign g10155 = (g3618&g1795);
assign g22493 = ((~g17042)&(~g21899));
assign II26532 = (g18561)|(g18514)|(g18458);
assign g29705 = ((~g6104)&(~g29583)&(~g25339));
assign g15675 = ((~II21926));
assign g16739 = ((~g14922));
assign g11808 = ((~g10996));
assign II16215 = ((~g3462));
assign II23682 = ((~g14966));
assign g26276 = ((~II34230));
assign g18429 = ((~g14831));
assign II24055 = ((~g14286))|((~II24053));
assign g13272 = ((~g10127));
assign II13987 = ((~g2451));
assign g26263 = (g4476&g25502);
assign II15392 = ((~g2556));
assign II31949 = ((~g23943));
assign g21982 = ((~II28541));
assign II17898 = ((~g6643));
assign g5638 = ((~II14094));
assign II25700 = ((~g1435))|((~g18297));
assign II15490 = ((~g3251));
assign II39886 = ((~g30284));
assign g28213 = ((~II36888));
assign g25356 = (g5898&g24607);
assign g22500 = ((~II29046));
assign g20440 = ((~II26871));
assign g27711 = ((~II36144));
assign g16997 = (g7578&g15352);
assign g22658 = ((~II29280));
assign g20655 = ((~II27246));
assign g10662 = (g3678&g5306);
assign g25267 = ((~g24884)&(~g17936));
assign g20391 = ((~g17537));
assign g18851 = ((~g15317));
assign g16346 = (g295&g11972);
assign g10849 = ((~II17698));
assign g21533 = (g17724&g18179&g19799&II28068);
assign g21197 = (g5912&g19330);
assign g27793 = ((~II36240));
assign g18901 = ((~g15499));
assign g30254 = ((~g16242)&(~g30088));
assign g21091 = (g20250&g12166);
assign g21498 = ((~II28038));
assign II29475 = ((~g21005));
assign g21989 = ((~g21048))|((~g18623));
assign g15022 = ((~g11781));
assign g24873 = ((~II32560))|((~II32561));
assign II29942 = ((~g22548));
assign II25741 = ((~g1439))|((~II25740));
assign g5881 = ((~g2378));
assign g7963 = ((~II15271));
assign g14332 = ((~g12068));
assign g30732 = ((~II40484));
assign g22308 = ((~g20182)&(~g21812));
assign g12546 = ((~g8693));
assign g8304 = ((~g3773));
assign g19333 = (g16954)|(g16602)|(g16560);
assign g25518 = (g24489&g20447);
assign II34990 = ((~g26573));
assign g25068 = ((~g23803))|((~g5556));
assign II30398 = ((~g22840));
assign g13541 = ((~g13274));
assign g8658 = ((~II15850));
assign g18858 = ((~g15346));
assign II14134 = ((~g1018));
assign g22118 = ((~g19521))|((~g21269))|((~g19542));
assign g30898 = ((~II40946));
assign II19813 = ((~g10649));
assign g3249 = ((~II13143));
assign II18587 = ((~g8718));
assign II14704 = ((~g2818));
assign g10506 = (g3494&g5047);
assign II40937 = ((~g30833));
assign g25911 = ((~g24962));
assign g16586 = ((~g14507));
assign g8431 = (g3254&g237);
assign g19189 = ((~II25412));
assign II31274 = ((~g22249));
assign g25054 = ((~g23955))|((~g6751));
assign g16607 = (g15022&g15096);
assign II40862 = ((~g30773));
assign g26354 = ((~II34313));
assign II16854 = ((~g7195));
assign g23712 = ((~II30878));
assign g22797 = ((~II29575));
assign g23639 = (g21825&g22805);
assign g30870 = ((~II40862));
assign II24641 = ((~g15210))|((~II24639));
assign g29777 = ((~g29478)&(~g29225));
assign g3994 = ((~g2848));
assign II31829 = ((~g23871));
assign II34162 = ((~g25684));
assign II31505 = ((~g23589));
assign g29772 = ((~g29473)&(~g29203));
assign II18780 = ((~g10870));
assign g30739 = ((~II40501));
assign g18969 = ((~II25015));
assign II41129 = ((~g30973));
assign g30250 = ((~g16163)&(~g30083));
assign g21055 = ((~g19904)&(~g18129));
assign g24849 = ((~g24254))|((~g24257));
assign g5889 = ((~II14343));
assign g15404 = ((~II21666));
assign II28206 = ((~g20067));
assign g12711 = ((~II19803));
assign g23128 = (g5943&g21079);
assign g23116 = ((~II29863));
assign g12013 = ((~g10772));
assign g22044 = ((~g21311)&(~g19571));
assign II31673 = ((~g23492));
assign II30493 = ((~g23030));
assign II37842 = ((~g28501));
assign g20123 = (g18478)|(g18395)|(II26571);
assign g27926 = (g13992&g27428);
assign g30128 = (g30062&g20722);
assign g14551 = ((~g12215));
assign g6898 = ((~g2993));
assign g10224 = (g6783&g4538);
assign g6441 = ((~g2366));
assign II33485 = ((~g25034));
assign g11744 = ((~g9241)&(~g9301)&(~g9364));
assign g13250 = ((~g10021));
assign II39240 = ((~g29691));
assign g5945 = ((~g2190));
assign g18764 = ((~g15055));
assign g26073 = ((~g25438))|((~g25405))|((~g25291));
assign g12776 = ((~g10766));
assign g13345 = (g5746&g11324);
assign g23855 = (g22954&g9767);
assign II37238 = ((~g28179));
assign g12288 = ((~g10569)&(~g10614)&(~g10651));
assign g20211 = (g13714&g13791&II26645);
assign g28717 = (g28461&g19346);
assign II22044 = ((~g11733));
assign g4973 = ((~g2108));
assign II36042 = ((~g26960));
assign II34836 = ((~g26480));
assign g28497 = (g18573&g28190);
assign g24366 = ((~II31772));
assign g11499 = ((~II18473));
assign g29995 = (g29893&g8434);
assign g13205 = ((~g9641));
assign g19777 = (g17927&g16056);
assign g5431 = ((~g3211));
assign g29445 = ((~II38716));
assign g22270 = (g92&g21529);
assign g20763 = ((~II27352));
assign g4405 = ((~g1801));
assign II19119 = ((~g9202));
assign II31595 = ((~g23561));
assign II20310 = ((~g9067));
assign II24520 = ((~g6435))|((~g14234));
assign g23293 = ((~II30332));
assign g29013 = ((~g28671)&(~g11607));
assign g26565 = ((~g25536));
assign g19873 = (g1365&g18929);
assign II25768 = ((~g17139));
assign g28688 = ((~II37611));
assign g12916 = (II19971&II19972);
assign gbuf109 = (g1254);
assign g29713 = ((~g6104)&(~g29583)&(~g25332));
assign II29451 = ((~g20997));
assign g4779 = ((~g1211));
assign g16337 = ((~g12328));
assign g16554 = ((~g14395));
assign g28238 = ((~II36963));
assign II37502 = ((~g27768));
assign g12234 = ((~g10479)&(~g10540)&(~g10599));
assign II36560 = ((~g27285));
assign g7518 = ((~g2354));
assign g19862 = (g2746&g18925);
assign g30886 = ((~II40910));
assign g29149 = ((~II38190));
assign g19219 = ((~g18165)&(~g15753));
assign g4020 = ((~g700));
assign g25885 = ((~g4809)&(~g14985)&(~g25091));
assign g17537 = ((~II23625));
assign g22237 = ((~g20644));
assign g11544 = ((~II18608));
assign II36510 = ((~g27271));
assign g10598 = (g7426&g5224);
assign g28813 = ((~g28497)&(~g28066));
assign g30553 = ((~II40239));
assign g21381 = (g15022&g20381);
assign g23744 = ((~II30938));
assign g28002 = ((~g26032)&(~g27246));
assign g21342 = (g9488&g20342);
assign II40604 = ((~g30614))|((~II40603));
assign g23737 = ((~II30925));
assign g30896 = ((~II40940));
assign g30278 = ((~g16420)&(~g30112));
assign II33440 = ((~g25048));
assign g19141 = ((~g3088))|((~g16825));
assign g19639 = (g4061&g17416);
assign g7142 = ((~g8));
assign g7973 = ((~g3068));
assign g22672 = ((~II29310));
assign g14352 = ((~g12081));
assign g30914 = ((~II40994));
assign g19504 = ((~g16785));
assign g10385 = (g7162&g4800);
assign g4731 = ((~g2782));
assign II23192 = ((~g13999))|((~II23190));
assign g29806 = ((~II39270));
assign g30404 = ((~g30006)&(~g30132));
assign g6083 = ((~II14596));
assign g12530 = ((~g8667));
assign g20626 = ((~II27203));
assign II15896 = ((~g3878));
assign II21534 = ((~g13045));
assign g27404 = ((~II35744));
assign II36945 = ((~g27793));
assign g19717 = (g2072&g18847);
assign g25454 = ((~II33278));
assign II21354 = ((~g11798));
assign g22679 = (g14107&g21541);
assign g10961 = ((~g5978));
assign II35780 = ((~g27124));
assign g18466 = ((~II24507));
assign II16763 = ((~g6945));
assign g28089 = ((~II36702));
assign g7488 = ((~II15015));
assign II36542 = ((~g27280));
assign g30449 = (g30159&g11151);
assign g25496 = ((~II33324));
assign g16971 = ((~II22912));
assign g29944 = (g29782&g28889);
assign g25628 = (g21008&g25115);
assign g5030 = ((~g586));
assign II17825 = ((~g7483));
assign g11170 = ((~II18088));
assign g28796 = ((~II37757));
assign g12965 = ((~g9006));
assign II34749 = ((~g26205));
assign g14976 = ((~g12248));
assign g14478 = ((~g12162));
assign g8897 = ((~II16169));
assign g28231 = ((~II36942));
assign g12343 = ((~II19510));
assign g17653 = (g4483&g15329);
assign g10008 = (g6232&g4208);
assign II33463 = ((~g25030));
assign II27375 = ((~g19431));
assign II16098 = ((~g6084));
assign g15996 = ((~g12955))|((~g7358));
assign gbuf102 = (g1199);
assign II29600 = ((~g21720));
assign g11696 = ((~g9534))|((~g3366));
assign II40453 = ((~g30600));
assign g30435 = ((~II39985));
assign g14904 = ((~g11870));
assign g13023 = (g8027&g10482);
assign g18374 = ((~g14385));
assign g23618 = (g22608&g20383);
assign g22203 = ((~II28754))|((~II28755));
assign g25028 = ((~g23644))|((~g5438));
assign g8836 = ((~II16068));
assign g10604 = (g3338&g620);
assign g4194 = ((~g2249));
assign g16180 = ((~g12904));
assign g5865 = ((~g1466));
assign II18034 = ((~g6838));
assign g18013 = (g5064&g15612);
assign g13485 = (g6022&g12211);
assign g17000 = ((~II22963))|((~II22964));
assign g27346 = ((~g27105)&(~g26488));
assign g27603 = ((~g27179)&(~g17031));
assign g11020 = ((~g6029));
assign II32500 = ((~g24069))|((~II32498));
assign g30903 = ((~II40961));
assign g29427 = ((~II38662));
assign II27035 = ((~g19556));
assign g24277 = ((~II31505));
assign g26784 = (g24941&g26521&g13637);
assign g10526 = (g7358&g5101);
assign g6980 = ((~II14877));
assign g27123 = ((~g26583)&(~g17031));
assign g25260 = ((~g24858)&(~g17737));
assign g29440 = ((~II38701));
assign g13504 = (g6038&g12266);
assign gbuf138 = (g1738);
assign g16126 = ((~g12854));
assign II35467 = ((~g26834));
assign g18353 = ((~g13918));
assign g13321 = ((~II20386));
assign II38510 = ((~g28778));
assign g26698 = ((~II34701));
assign II38223 = ((~g29106));
assign g18450 = ((~II24481));
assign g14402 = ((~g12108));
assign II14017 = ((~g1657));
assign II26494 = ((~g18102));
assign II19905 = ((~g8726));
assign g17968 = ((~II24006))|((~II24007));
assign II35711 = ((~g26974));
assign g17333 = ((~II23421));
assign g28698 = ((~II37641));
assign g22842 = (g3032&g21682);
assign g28304 = ((~II37161));
assign g22626 = ((~II29220));
assign g27190 = ((~II35407));
assign II20852 = ((~g12457));
assign g22801 = ((~II29585));
assign g16383 = (g5928&g12023);
assign g7345 = ((~g3139));
assign II25150 = ((~g18991));
assign g6082 = ((~II14593));
assign g30959 = ((~g30923)&(~g30949));
assign II23257 = ((~g9795))|((~II23256));
assign II32556 = ((~g23329));
assign g26056 = ((~II33954));
assign g30122 = ((~II39631));
assign g6672 = ((~g464));
assign II18247 = ((~g6945));
assign g29256 = (g28859&g8894);
assign II19611 = ((~g9276));
assign II28978 = ((~g21740));
assign g23914 = (g22975&g10087);
assign g29198 = ((~g15047)&(~g28898));
assign g8394 = (g3410&g906);
assign g26110 = ((~g6068)&(~g24183)&(~g25305));
assign g7915 = ((~g2704));
assign g19033 = ((~II25162));
assign g12742 = ((~g8813));
assign g22444 = ((~II28988));
assign g30985 = ((~II41129));
assign g21857 = ((~g18079))|((~g19192))|((~g19200));
assign II36789 = ((~g27344));
assign II29046 = ((~g21776));
assign g8224 = ((~g1523));
assign II24717 = ((~g14497))|((~II24716));
assign II31141 = ((~g22777));
assign g29333 = ((~g28719)&(~g19131));
assign g24177 = ((~g22603));
assign II40793 = ((~g30821));
assign g11135 = ((~II18049));
assign g21622 = (g16520&g19505&g14186);
assign II25660 = ((~g17204));
assign g25487 = (g24485&g20425);
assign g11095 = ((~II18007));
assign g4338 = ((~II13430));
assign g30666 = ((~g16369)&(~g30476));
assign g12532 = ((~g8670));
assign II13433 = ((~g105));
assign g20480 = (g17313&g11827);
assign g10370 = (g3366&g4763);
assign g11917 = ((~g9957)&(~g10080)&(~g10171));
assign g28341 = ((~II37228));
assign II31934 = ((~g24068));
assign g24717 = ((~g23886)&(~g22754));
assign g13119 = ((~g9822))|((~g7358));
assign II29897 = ((~g23116));
assign g19177 = ((~g17713)&(~g15442));
assign g25063 = ((~g24014))|((~g7391));
assign g5831 = ((~g1887));
assign g14007 = (g7673&g12915);
assign g23717 = (g22680&g20433);
assign g9277 = ((~g5995));
assign II35064 = ((~g26531));
assign g11508 = ((~II18500));
assign g21217 = ((~g19125));
assign g19301 = ((~g16622));
assign II26429 = (g17979)|(g17887)|(g17807);
assign II35500 = ((~g26890));
assign g30578 = ((~II40288));
assign g15441 = ((~g12418));
assign g18795 = ((~g15151));
assign g19549 = (g7950&g17230);
assign g28635 = ((~g28189)&(~g17031));
assign g18855 = ((~g15332));
assign g16578 = ((~g14478));
assign g30261 = ((~g16342)&(~g30095));
assign g8253 = ((~g3053));
assign g26557 = ((~g13818)&(~g25286));
assign g22145 = ((~g21411)&(~g19736));
assign II28272 = ((~g14431))|((~II28271));
assign II41024 = ((~g30765));
assign g27060 = (g22016&g26626);
assign II31766 = ((~g23792));
assign g26011 = ((~II33885));
assign g29481 = (g21508&g29283);
assign II23830 = ((~g13558));
assign g12315 = ((~II19482));
assign g20503 = (g17507&g13817);
assign g22028 = ((~g21291)&(~g19554));
assign gbuf68 = (g520);
assign g23533 = ((~g22939))|((~g14618))|((~g10754));
assign g13454 = ((~II20661));
assign II36271 = ((~g27549))|((~II36270));
assign g9286 = ((~g6197));
assign g28245 = ((~II36984));
assign g10868 = ((~II17721));
assign g30667 = ((~g16370)&(~g30477));
assign II27739 = (g19379&g19348&g19325);
assign g25256 = ((~g24840)&(~g23721));
assign II30095 = ((~g22733));
assign g9078 = (g3462&g7652);
assign g21350 = (g9203&g20348);
assign g24324 = ((~II31646));
assign II32432 = ((~g24052))|((~II32430));
assign g4743 = ((~g575));
assign II23839 = ((~g14985));
assign g20363 = ((~g17436));
assign g8452 = ((~II15654));
assign g19346 = ((~g16644));
assign g24571 = (g18630&g23435&g20005);
assign g23023 = ((~g14256)&(~g14175)&(~g21123));
assign II17297 = ((~g6130));
assign g22709 = ((~II29383));
assign II40940 = ((~g30828));
assign II29052 = ((~g21780));
assign II30326 = ((~g22774));
assign g9520 = (g6232&g8197);
assign g18754 = ((~g13655)&(~g11816));
assign g10013 = (g3306&g4221);
assign g14626 = ((~g12306));
assign g30523 = ((~II40149));
assign II20664 = ((~g13325));
assign g25014 = ((~g23694))|((~g5473));
assign g14438 = ((~g12124));
assign g10324 = (g6838&g4708);
assign II16306 = ((~g7015));
assign g15360 = ((~II21629));
assign g25582 = ((~II33405));
assign II39835 = ((~g30271));
assign g16160 = (g8286&g11836);
assign g30088 = (g29844&g11138);
assign II26182 = ((~g18308));
assign II40573 = ((~g30632))|((~II40571));
assign g12354 = ((~g8381));
assign II39234 = ((~g29689));
assign g29439 = ((~II38698));
assign gbuf135 = (g1723);
assign II34091 = ((~g25217));
assign II29265 = ((~g20927));
assign g18200 = ((~g14183));
assign g18895 = ((~II24923));
assign g12892 = ((~g8928));
assign II17599 = (g7566&g7583&g7587);
assign g25825 = ((~g24619));
assign g30872 = ((~II40868));
assign g30340 = (g30207&g8372);
assign II31181 = ((~g22200));
assign g23107 = (g21813)|(g21807);
assign g12082 = ((~g10290)&(~g10368)&(~g10435));
assign g28278 = ((~II37083));
assign g20095 = ((~g16507)&(~g16895));
assign g30967 = ((~g30954));
assign g8872 = ((~II16134));
assign g15754 = (g7837&g13308);
assign II16735 = (g5856&g4338&g4339&g5141);
assign g26464 = (g5238&g25821);
assign g23727 = ((~II30905));
assign g13081 = ((~g9968))|((~g7488));
assign II14612 = ((~g1779));
assign II23729 = ((~g14337));
assign g19355 = (g17136&g8605);
assign g25248 = ((~g24818)&(~g23664));
assign g29816 = (g29759&g13883);
assign g12279 = ((~II19449));
assign g12033 = ((~g10199)&(~g10284)&(~g10362));
assign g17645 = ((~II23729));
assign g17989 = (g5035&g15596);
assign g5173 = ((~g1829));
assign g29922 = ((~g29744)&(~g22367));
assign g25606 = ((~II33431));
assign g29987 = (g29889&g8369);
assign g20421 = ((~g17649));
assign II25144 = ((~g18984));
assign II17692 = ((~g8107));
assign g10391 = (g3618&g1816);
assign g9227 = ((~g5587));
assign g28937 = ((~II37906));
assign g27275 = ((~g27003)&(~g26310));
assign g26422 = (g5104&g25746);
assign g13442 = ((~II20625));
assign II40688 = ((~g30644));
assign g11132 = ((~II18046));
assign II21262 = ((~g11713));
assign g18689 = (g14922&g13724&g13764&g16360);
assign g30053 = ((~g29963)&(~g16286));
assign II22578 = ((~g14746));
assign g13319 = ((~II20382));
assign g8869 = (g6776&g5552);
assign II27549 = ((~g20353));
assign g24292 = ((~II31550));
assign g21341 = (g9613&g20341);
assign II39142 = ((~g29581));
assign g26223 = ((~II34159));
assign g4202 = ((~g42));
assign g17496 = ((~II23584));
assign II38863 = ((~g29178));
assign II33003 = ((~g24956));
assign g24771 = ((~II32296))|((~II32297));
assign g10064 = (g7015&g1792);
assign g29229 = (g9293&g28791);
assign g9892 = (g3306&g414);
assign g26744 = ((~II34839));
assign II31472 = ((~g23548));
assign g23669 = ((~II30813));
assign II24030 = ((~g14086))|((~II24028));
assign g16520 = ((~g14273)&(~g14459));
assign g22986 = ((~g21382));
assign g22920 = ((~g21869))|((~g21864))|((~g21888));
assign II20628 = ((~g13394));
assign g15806 = ((~g12565))|((~g6314));
assign g25767 = ((~II33600));
assign g15151 = ((~g12005));
assign II35906 = ((~g14831))|((~II35904));
assign g19953 = (g7566&g18334);
assign g6221 = ((~g2628));
assign g27311 = ((~g27053)&(~g26396));
assign g19739 = (g4369&g17588);
assign g27168 = ((~II35373));
assign g12247 = ((~g10499)&(~g10559)&(~g10605));
assign g28333 = (g27882&g20772);
assign g21161 = (g20212&g12343);
assign g8724 = (g3650&g7862);
assign g30564 = ((~II40272));
assign g25352 = ((~g24875));
assign g12094 = ((~II19274));
assign g15606 = ((~II21862));
assign g8344 = ((~II15546));
assign II38217 = ((~g29105));
assign g5122 = ((~g2670));
assign g25899 = ((~g24928));
assign II16273 = ((~g3618));
assign II33424 = ((~g25023));
assign g11056 = ((~II17975));
assign g12149 = ((~g8336));
assign g30726 = ((~II40468));
assign g10423 = (g5438&g4885);
assign II22953 = ((~g15210))|((~II22952));
assign g29976 = ((~II39466));
assign g13265 = ((~g8568));
assign II35533 = ((~g26921));
assign II34051 = ((~g25204));
assign II29987 = ((~g22703));
assign g16572 = ((~II22640));
assign g27678 = ((~g26800)&(~g10133));
assign g29623 = ((~g14130)&(~g29264));
assign g23542 = ((~II30586));
assign g6068 = ((~g499));
assign g19563 = ((~II25994));
assign g26680 = ((~II34647));
assign II40892 = ((~g30831));
assign g20972 = ((~g19774)&(~g17752));
assign g8156 = ((~g1867));
assign g5678 = (g325&g379);
assign II19429 = ((~g10617));
assign g17973 = (g11623)|(g15659);
assign g17594 = ((~II23682));
assign II31487 = ((~g23557));
assign g30900 = ((~II40952));
assign g18383 = ((~II24400))|((~II24401));
assign g18207 = ((~g14207));
assign II24273 = ((~g13922))|((~II24271));
assign g19618 = (g3972&g17369);
assign g10584 = (g7053&g1985);
assign g21184 = ((~II27749));
assign g13872 = ((~g11780));
assign II36075 = ((~g27494));
assign II38235 = ((~g29118));
assign g12984 = (g9968)|(g3866);
assign II40727 = ((~g30657));
assign II40859 = ((~g30770));
assign g26764 = (g16632&g26525&g13649);
assign g13056 = (g4092&g10646);
assign g3242 = ((~II13122));
assign g28463 = (g28137&g9401);
assign II36551 = ((~g27282));
assign II32608 = ((~g18038))|((~II32607));
assign g23472 = ((~II30516));
assign II36347 = ((~g27630));
assign g25058 = ((~g23984))|((~g7053));
assign II14030 = ((~g182));
assign g27478 = ((~g26754)&(~g24432));
assign II20451 = ((~g10908));
assign II24373 = ((~g14454))|((~II24372));
assign II24453 = ((~g6142))|((~II24452));
assign g6574 = ((~II14786));
assign g5801 = ((~II14249));
assign g28851 = (g27892&g28618);
assign g9523 = (g6232&g8206);
assign g8952 = ((~II16258));
assign II14306 = ((~g97));
assign g18932 = ((~II24966));
assign g22102 = ((~g21362)&(~g19655));
assign g6040 = ((~II14513));
assign II36724 = ((~g27329));
assign g23549 = ((~II30601));
assign g11782 = ((~g10963));
assign g21174 = (g20223&g12363);
assign g4517 = ((~g1390));
assign g15949 = ((~g12711))|((~g6838));
assign g19738 = (g4366&g17585);
assign g28616 = ((~g27847));
assign g20914 = ((~g19673)&(~g17541));
assign II24290 = ((~g13895))|((~g9203));
assign II40745 = ((~g30663));
assign g21722 = ((~g20198))|((~g6519));
assign g28646 = ((~g27956));
assign g13764 = ((~g12461));
assign g19411 = ((~II25830))|((~II25831));
assign g18106 = (g5164&g15672);
assign g4322 = ((~g2839));
assign II28497 = ((~g21399));
assign II25819 = ((~g1448))|((~g18509));
assign g19913 = (g18247&g16236);
assign II30197 = ((~g22716));
assign g23898 = (g18390&g23075);
assign g27998 = ((~II36483));
assign g26966 = (g13963&g26196);
assign g9106 = (g7015&g7715);
assign II33265 = ((~g24925));
assign II33316 = ((~g24434));
assign g12027 = ((~II19208));
assign II35369 = ((~g26144));
assign g22805 = ((~g21894));
assign g29383 = ((~g28998));
assign II29556 = ((~g21033));
assign g23494 = (g18328&g22721);
assign g27008 = (g22050&g26581);
assign g27396 = (g692&g27135);
assign g5511 = ((~II14017));
assign g23775 = ((~II30979));
assign g23256 = ((~II30221));
assign g21818 = (g16736&g19641&g14863);
assign II23028 = ((~g15366))|((~II23027));
assign II28003 = ((~g19957));
assign g13549 = ((~g12611))|((~g3410));
assign g23227 = ((~II30134));
assign g7742 = ((~g1783));
assign g8793 = ((~II15995));
assign g17166 = (g7721&g14214);
assign g30451 = (g30155&g11163);
assign g8574 = ((~g3866))|((~g3834));
assign g11787 = ((~g10969));
assign g25936 = ((~g25000))|((~g5556));
assign g25353 = ((~g24904));
assign g20986 = ((~II27537));
assign g18053 = ((~II24077))|((~II24078));
assign II30716 = ((~g22061));
assign g24637 = ((~g23665)&(~g22587));
assign II16238 = ((~g7936));
assign g10298 = (g3462&g1122);
assign g29796 = ((~II39240));
assign g15095 = ((~II21420));
assign g22127 = ((~g21390)&(~g19702));
assign g8438 = (g6519&g921);
assign g23220 = ((~II30113));
assign II29090 = ((~g21772));
assign g17243 = ((~II23329));
assign g23968 = ((~g22852))|((~g13978));
assign g21540 = (g20542)|(g16895)|(g14186);
assign II34647 = ((~g26164));
assign II23769 = ((~g15899));
assign g23320 = ((~g23066))|((~g23051));
assign II23114 = ((~g9356))|((~II23113));
assign g28468 = (g18265&g28172);
assign II30263 = ((~g22768));
assign gbuf127 = (g1833);
assign II18289 = ((~g8102))|((~II18287));
assign g21635 = (g7549&g20496);
assign g11569 = ((~II18683));
assign g23154 = ((~II29915));
assign g11562 = ((~II18662));
assign II37712 = ((~g28512));
assign II13977 = ((~g2436));
assign g12844 = ((~II19905));
assign II30713 = ((~g22060));
assign g20124 = ((~II26574));
assign II20844 = ((~g12524));
assign g19264 = (g17830)|(g17919);
assign g22401 = ((~g21533));
assign g19713 = (g4272&g17537);
assign g12201 = ((~II19377));
assign II26947 = ((~g17429));
assign g30673 = ((~g16402)&(~g30490));
assign g24424 = ((~II31946));
assign g23641 = ((~II30779));
assign g29676 = ((~g29540)&(~g29320));
assign g5428 = ((~g3210));
assign g6911 = ((~II14857));
assign g14829 = ((~II21326));
assign II34725 = ((~g26239));
assign II15620 = ((~g3722));
assign g11836 = ((~g11042));
assign g19895 = (g686&g18945);
assign II36032 = ((~g27113));
assign g11848 = ((~II19030));
assign g5715 = ((~g541));
assign g14559 = ((~g13002));
assign g24210 = ((~g22696));
assign g7083 = ((~g1664));
assign g7899 = ((~g3066));
assign g14837 = ((~g12145));
assign g12388 = ((~g10709)&(~g10727)&(~g10745));
assign g19294 = (g16895)|(g16546)|(g16507);
assign g27112 = (g22157&g26662);
assign II32345 = ((~g17815))|((~g24002));
assign g18431 = ((~II24453))|((~II24454));
assign II34854 = ((~g26507));
assign g17633 = (g4444&g15314);
assign g24038 = ((~g4985)&(~g13602)&(~g23061));
assign g5654 = ((~g809));
assign II37626 = ((~g28393));
assign II13224 = ((~g2383));
assign g7336 = ((~g1476));
assign II26311 = (g18353&g13958&g14011);
assign g28126 = ((~II36803));
assign g7348 = ((~g451));
assign g17457 = ((~II23545));
assign g15293 = ((~II21569));
assign g19805 = (g17903&g16088);
assign II31011 = ((~g22151));
assign g21964 = ((~II28518));
assign g22614 = (g13963&g21477);
assign g26195 = ((~II34111));
assign II20676 = ((~g11616));
assign II26993 = ((~g19159));
assign g12974 = (II20021&II20022);
assign g19162 = ((~g17485)&(~g15243));
assign g9044 = ((~II16363));
assign g28438 = (g17882&g27919);
assign II30125 = ((~g22792));
assign gbuf152 = (g1903);
assign g11528 = ((~II18560));
assign g20512 = (g17445&g13836);
assign II26334 = ((~g18977));
assign g25171 = ((~II32991));
assign g12473 = ((~g8580));
assign g13790 = (g7475&g12558);
assign g8775 = ((~II15971));
assign g13037 = ((~g9676))|((~g6980));
assign g21774 = (g19121)|(g16884)|(g14776);
assign g11760 = ((~g9319)&(~g9382)&(~g9461));
assign g21873 = ((~g18395))|((~g19227))|((~g19234));
assign II32284 = ((~g17815))|((~g23953));
assign g13633 = ((~g12984))|((~g3834));
assign II23326 = ((~g15758));
assign II37158 = ((~g28110));
assign g22622 = ((~II29212));
assign II17828 = ((~g7389));
assign g16421 = (g5962&g12087);
assign g30776 = ((~II40594));
assign II25588 = (g17201)|(g17192)|(g17180);
assign g21036 = ((~II27593));
assign g23166 = ((~II29951));
assign g11606 = ((~II18780));
assign g30462 = (g30171&g11237);
assign g12176 = ((~g8372));
assign g24244 = (g14144)|(g22317);
assign g21677 = ((~g20099)&(~g14309)&(~g14402));
assign g26126 = ((~g6068)&(~g24183)&(~g25368));
assign gbuf146 = (g1778);
assign II27173 = ((~g20440));
assign g14214 = ((~II21119));
assign II36213 = ((~g27571));
assign g25394 = ((~g24753));
assign II26354 = (g18388&g18312&g18224);
assign g17300 = ((~II23386));
assign g11189 = ((~II18114))|((~II18115));
assign g18319 = ((~II24326))|((~II24327));
assign II35957 = ((~g26947));
assign g12089 = ((~g11441));
assign II31000 = ((~g22847));
assign g28225 = ((~II36924));
assign g16529 = ((~g14301));
assign II36951 = ((~g27992));
assign g7901 = ((~II15222));
assign g4346 = ((~g432));
assign II19771 = ((~g10038));
assign g12482 = ((~g9057)&(~g9073)&(~g9082));
assign g16048 = (g6170&g11762);
assign g19092 = (g14776&g18670&g18692&g16293);
assign II23125 = ((~g13866))|((~II23123));
assign II20320 = ((~g10792));
assign g16416 = (g5957&g12078);
assign II23142 = ((~g9407))|((~g13991));
assign g8407 = (g6574&g1603);
assign II39261 = ((~g29697));
assign g11663 = ((~g9095)&(~g9104)&(~g9112));
assign II31823 = ((~g23870));
assign g28728 = ((~g28422)&(~g27904));
assign II16832 = ((~g6081));
assign g26243 = (g4372&g25484);
assign g30934 = ((~g30759)&(~g30761));
assign g13598 = ((~II20816));
assign II39044 = ((~g29511));
assign g26831 = ((~II34964));
assign II31805 = ((~g24248));
assign II23981 = ((~g14292))|((~g9216));
assign II28341 = (g19106)|(g19101)|(g19095);
assign g22232 = ((~II28800));
assign II36924 = ((~g28026));
assign II19573 = ((~g8835));
assign g24481 = ((~g23618)&(~g19696));
assign II40468 = ((~g30672));
assign II38502 = ((~g28773));
assign g20448 = ((~g17767));
assign g8366 = ((~II15568));
assign g15844 = ((~g12565))|((~g6232));
assign g9058 = ((~II16372));
assign II39136 = ((~g29611));
assign g8056 = ((~g146));
assign g17081 = (g7614&g15578);
assign g27798 = ((~g27632)&(~g1223));
assign II30008 = ((~g22785));
assign g17310 = ((~II23398));
assign g29401 = ((~II38594));
assign g16142 = ((~g13057));
assign g22573 = ((~II29135));
assign g24528 = ((~g23851)&(~g22722));
assign g24755 = (g9569&g24108);
assign II40769 = ((~g30803));
assign II23386 = ((~g13469));
assign g25178 = (g24623&g20634);
assign g17514 = ((~II23602));
assign g29472 = (g21461&g29268);
assign g11986 = ((~g11294));
assign g27227 = ((~II35518));
assign II29996 = ((~g22729));
assign g23157 = ((~II29924));
assign g17624 = ((~II23712));
assign II15472 = ((~g3245));
assign g26159 = ((~II34051));
assign g23095 = ((~g21671));
assign g6052 = ((~II14535));
assign II40594 = ((~g30705));
assign g28945 = ((~II37912));
assign g11590 = ((~II18746));
assign g16489 = ((~II22569));
assign g24140 = ((~g22494));
assign g25371 = (g5937&g24619);
assign g30751 = ((~II40531));
assign g29766 = ((~g29467)&(~g19142));
assign g30945 = (g30931&g20754);
assign g8536 = (g6369&g891);
assign g29980 = (g29881&g8324);
assign g9763 = (g6314&g4012);
assign g10460 = (g3678&g4964);
assign II17822 = ((~g7478));
assign II40224 = ((~g30336));
assign g24834 = ((~g23455));
assign g24940 = ((~II32696))|((~II32697));
assign II24407 = ((~g6298))|((~g14119));
assign g16505 = (g14776&g14797&g16142&g16243);
assign II39948 = ((~g30303));
assign g28315 = ((~II37194));
assign g16428 = (g1676&g12105);
assign g30117 = (g29877&g11465);
assign g13957 = ((~g10730))|((~g12473));
assign II22679 = ((~g14669));
assign II14006 = ((~g963));
assign g10810 = ((~g5711)&(~g5758)&(~g5807));
assign g5799 = ((~II14243));
assign g23846 = ((~II31088));
assign g11713 = ((~g10481))|((~g9144));
assign II33897 = ((~g25851));
assign g13221 = ((~g9790));
assign II23380 = ((~g15809));
assign II14562 = ((~g398));
assign g19664 = (g4130&g17454);
assign g21303 = (g9595&g20292);
assign gbuf34 = (g286);
assign II17801 = ((~g8107));
assign II21083 = ((~g12535));
assign g27462 = ((~g26892)&(~g24622));
assign g24821 = (g9795&g24163);
assign g21505 = ((~II28043));
assign II21389 = ((~g12883));
assign g28326 = (g27865&g22274);
assign g29488 = (g21544&g29295);
assign g16474 = ((~II22524));
assign g24442 = ((~g23644))|((~g3306));
assign g24285 = ((~II31529));
assign g23066 = ((~g21138)&(~g19303)&(~g19320));
assign g11597 = ((~II18767));
assign II40760 = ((~g30722));
assign g11101 = ((~II18013));
assign g18505 = ((~II24560));
assign II24179 = ((~g13873))|((~II24178));
assign II30810 = ((~g22090));
assign g23851 = (g7329&g23048);
assign g29434 = ((~II38683));
assign g15726 = ((~II21974));
assign II27346 = ((~g19431));
assign g28262 = ((~II37035));
assign II19605 = ((~g10797));
assign g16590 = (g14936&g15003&g16325&g16404);
assign g27034 = (g22069&g26605);
assign g18970 = ((~II25018));
assign II28813 = ((~g21502));
assign g28426 = (g28128&g9170);
assign g21800 = (g18665)|(g20270)|(g20248)|(g18647);
assign g14090 = ((~g11939));
assign g29378 = ((~g28972));
assign II28518 = ((~g20985));
assign g19839 = (g666&g18909);
assign g8013 = ((~g1855));
assign g6289 = ((~g1228));
assign g28731 = ((~g28423)&(~g27908));
assign g22126 = ((~g21389)&(~g19701));
assign g9908 = (g3410&g4136);
assign g6895 = ((~II14848));
assign g23167 = ((~II29954));
assign g21024 = ((~II27577));
assign g25830 = ((~II33670));
assign g21204 = ((~g20123)&(~g20102));
assign g9931 = (g5512&g1789);
assign g25064 = ((~g23955))|((~g6751));
assign g23177 = ((~II29984));
assign g25763 = ((~II33596));
assign II16153 = ((~g3306));
assign g25853 = ((~g25081)&(~g21674));
assign g25444 = ((~g24641));
assign II29727 = ((~g20877));
assign g11948 = ((~g11231));
assign II18175 = ((~g7085));
assign g20402 = ((~g17573));
assign g24312 = ((~II31610));
assign II20351 = ((~g10804));
assign II21844 = ((~g13131));
assign gbuf213 = (g2623);
assign g26757 = ((~II34872));
assign g9664 = (g6519&g3960);
assign II40155 = ((~g30369));
assign g18718 = (g15003&g13774&g13805&g16404);
assign g16297 = ((~II22382));
assign II14182 = ((~g1712));
assign g5980 = ((~g201));
assign g19052 = ((~II25219));
assign II31781 = ((~g23838));
assign g19243 = (g16995)|(g16986)|(II25500);
assign g26167 = ((~II34063));
assign g23241 = ((~II30176));
assign gbuf120 = (g1520);
assign g13169 = ((~g9320));
assign g19067 = ((~g16554))|((~g16578));
assign g13581 = ((~II20805));
assign g10113 = (g6912&g4351);
assign g6059 = ((~II14556));
assign g27936 = (g4283&g27440);
assign gbuf181 = (g2361);
assign II16300 = ((~g3462));
assign g18728 = ((~g14910));
assign g19692 = (g4205&g17487);
assign II30544 = ((~g23092));
assign g15508 = (g5004&g13226);
assign g10205 = (g6678&g4492);
assign g12349 = ((~II19516));
assign g28035 = (g27599&g9916);
assign g11078 = ((~g6041));
assign g17896 = ((~g14352)&(~g16020));
assign g21253 = (g19608)|(g16728)|(g14811);
assign II16089 = ((~g6751));
assign g22634 = (g21939&g12765);
assign g11882 = ((~g9872)&(~g9956)&(~g10079));
assign g29517 = ((~II38881));
assign II24234 = ((~g14222))|((~g9613));
assign II27260 = ((~g19457));
assign g12088 = ((~g11438));
assign g20431 = ((~g17685));
assign II23131 = ((~g9391))|((~g13901));
assign g25295 = (g24704&g8780);
assign II25578 = ((~g780))|((~g18281));
assign II29415 = ((~g20981));
assign g27657 = (g27114&g11051);
assign II35905 = ((~g27051))|((~II35904));
assign II23243 = ((~g9737))|((~II23242));
assign II29625 = ((~g21056));
assign II23748 = ((~g14904));
assign II13190 = ((~g1236));
assign II18449 = ((~g10868));
assign g24506 = ((~g23776)&(~g22667));
assign II25623 = ((~g1466))|((~g18374));
assign g9760 = (g6314&g4003);
assign g17339 = (g8176&g15997);
assign g5754 = ((~g234));
assign g30809 = ((~II40679));
assign g24164 = ((~g22563));
assign II13203 = ((~g1689));
assign g28072 = ((~II36659));
assign g26750 = ((~II34857));
assign g15128 = ((~g12091));
assign II34146 = ((~g25232));
assign II22572 = ((~g15019));
assign g19824 = (g4714&g17785);
assign g10555 = (g3338&g5145);
assign g24145 = ((~g20956))|((~g22205));
assign g27142 = ((~g26254));
assign g24473 = ((~g23461)&(~g18407));
assign II14547 = ((~g384));
assign II29542 = ((~g21029));
assign II32943 = ((~g24583));
assign II13417 = ((~g2839));
assign II36568 = ((~g27287));
assign II13197 = ((~g1316));
assign g18951 = ((~g15691));
assign g18984 = ((~II25044));
assign g20369 = ((~g17465));
assign II31580 = ((~g23826));
assign g28013 = ((~II36516));
assign g25987 = ((~II33813));
assign g10368 = (g6912&g4757);
assign g13512 = ((~g12657))|((~g3566));
assign II19938 = (g9232&g9187&g9161&g9150);
assign g27528 = ((~II35905))|((~II35906));
assign II14660 = ((~g1211));
assign II24443 = ((~g14148))|((~g9507));
assign g29853 = ((~g29672));
assign II23055 = ((~g9264))|((~g13982));
assign g24553 = (g23429&g18007&g23071);
assign g5034 = ((~g614));
assign g16322 = (g5877&g11958);
assign g22206 = (g21895&g11976);
assign g10283 = (g3338&g573);
assign g4498 = ((~g817));
assign g15355 = ((~g12388));
assign g11348 = ((~II18302));
assign II19645 = ((~g10818));
assign g25102 = (g23444&g10915);
assign II18106 = ((~g7875))|((~g7855));
assign II26112 = ((~g16844));
assign II23226 = ((~g9649))|((~II23225));
assign g10109 = ((~II17081));
assign g30641 = ((~g16188)&(~g30438));
assign g11042 = ((~II17957));
assign g28414 = ((~g27748)&(~g22344));
assign g26380 = (g4948&g25672);
assign g4794 = ((~g1403));
assign g8637 = ((~II15827));
assign g4191 = ((~g2244));
assign g19416 = ((~II25847))|((~II25848));
assign g30648 = ((~g16252)&(~g30448));
assign g30282 = ((~g16430)&(~g30117));
assign g11555 = ((~II18641));
assign g24922 = (g2740&g23901);
assign g10161 = ((~II17125));
assign II34150 = ((~g25233));
assign gbuf85 = (g977);
assign g22870 = ((~g21293)&(~g20866));
assign g30292 = ((~g13477)&(~g29988));
assign g27339 = ((~g27093)&(~g26464));
assign g27174 = ((~g23494)&(~g26080));
assign II31862 = ((~g23718));
assign II17066 = ((~g3900));
assign g15020 = (g8090&g12561);
assign II18288 = ((~g8256))|((~II18287));
assign g29169 = ((~g28843)&(~g28398));
assign g10337 = ((~II17303));
assign g23106 = (g5857&g21050);
assign g25887 = ((~g4809)&(~g25091)&(~g18566)&(~g16164));
assign II31886 = ((~g23800));
assign g19020 = ((~II25123));
assign II20483 = ((~g9050));
assign g23513 = ((~g22911)&(~g5631));
assign II39332 = ((~g29705))|((~II39331));
assign g24252 = (g14259)|(g22342);
assign g27232 = ((~II35533));
assign II30305 = ((~g22746));
assign g5598 = ((~II14056));
assign g26063 = ((~II33961));
assign g15628 = ((~II21881));
assign II18835 = ((~g10834));
assign g4691 = ((~g1813));
assign g19847 = (g1352&g18915);
assign II40865 = ((~g30776));
assign II24215 = ((~g9711))|((~II24213));
assign g24532 = ((~g15545)&(~g23889));
assign II15642 = ((~g3566));
assign II25426 = ((~g18836));
assign II15935 = ((~g3878));
assign g15306 = ((~g12225));
assign g15560 = ((~g12343));
assign II34833 = ((~g26428));
assign II16587 = ((~g3462));
assign g29668 = ((~g29569));
assign g14691 = ((~II21267));
assign g25429 = ((~g24482)&(~g22319));
assign II21246 = ((~g11624));
assign g30843 = ((~II40781));
assign g5591 = ((~g3173));
assign II24028 = ((~g6201))|((~g14086));
assign g14541 = ((~g13001));
assign II23335 = ((~g16412));
assign g19285 = (g16749&g7642);
assign II34456 = ((~g25934));
assign II16601 = ((~g7015));
assign g12003 = ((~g11321));
assign g6442 = ((~II14755));
assign g27981 = ((~II36454));
assign II32560 = ((~g17927))|((~II32559));
assign II24709 = ((~g14502))|((~g15296));
assign g10643 = (g7488&g5283);
assign g7466 = ((~g3010));
assign II28080 = ((~g20487));
assign g20114 = (g17969&g9755);
assign II19800 = ((~g10574));
assign II14243 = ((~g3221));
assign gbuf61 = (g474);
assign g13096 = ((~g9968))|((~g7426));
assign g13648 = (g6294&g12513);
assign g22838 = ((~II29635));
assign g12420 = ((~g10986));
assign g25941 = ((~g24529)&(~g24540));
assign g29027 = ((~II37986));
assign g11085 = ((~II17995));
assign II40140 = ((~g30328));
assign g21864 = ((~g18147))|((~g19206))|((~g19215));
assign g24159 = ((~g22537));
assign g19741 = (g1339&g18856);
assign g10070 = ((~II17030));
assign g17798 = (g4591&g16099);
assign II28765 = ((~g21901))|((~g13552));
assign g26002 = ((~II33858));
assign g19008 = ((~II25089));
assign g12545 = ((~g8690));
assign g14071 = ((~g11934));
assign g24576 = ((~II32126));
assign II36545 = ((~g27281));
assign g18295 = ((~g14374));
assign g28689 = ((~II37614));
assign g26813 = ((~g15337)&(~g26302));
assign II29827 = ((~g21502));
assign g9301 = (g6314&g7990);
assign II13155 = ((~g51));
assign g30942 = ((~II41050));
assign g21155 = (g20140&g12336);
assign g13331 = ((~g8183)&(~g11332)&(~g11190)&(~g11069));
assign g18915 = ((~g15550));
assign g24798 = (g9649&g24148);
assign g18959 = ((~II25001));
assign g28750 = ((~g28436)&(~g27926));
assign g27332 = ((~g27084)&(~g26446));
assign g26525 = ((~g25340));
assign II27161 = ((~g20377));
assign g12502 = ((~g8640));
assign g21763 = ((~g20526)&(~g18503));
assign g10327 = (g5556&g4717);
assign g9440 = (g6232&g8129);
assign g21241 = ((~g19945));
assign II18359 = ((~g6838));
assign g15760 = ((~g12611))|((~g6369));
assign g30693 = ((~g13503)&(~g30364));
assign g22082 = ((~II28628));
assign g25998 = ((~II33846));
assign g26987 = ((~g26056));
assign g21230 = ((~g19266)&(~g19256));
assign g5606 = ((~g79));
assign II23162 = ((~g9453))|((~II23161));
assign g16705 = ((~g14849)&(~g14976));
assign g26353 = (g25923&g9752);
assign g22273 = (g21690&g12285);
assign g23036 = ((~g21558));
assign II23651 = ((~g13538));
assign g5927 = ((~g264));
assign g6750 = ((~II14822));
assign g8493 = (g6574&g1630);
assign g25620 = ((~II33445));
assign g29695 = ((~II39139));
assign g17183 = ((~g14132))|((~g14060));
assign g12523 = ((~g8296))|((~g7015));
assign g7013 = ((~g968));
assign g16357 = (g5907&g11994);
assign gbuf147 = (g1706);
assign g10041 = (g6369&g4234);
assign g23213 = ((~II30092));
assign II32468 = ((~g17903))|((~g24058));
assign g30531 = ((~II40173));
assign g14450 = ((~g12146));
assign g21917 = ((~II28435));
assign II37765 = ((~g28512));
assign g28170 = ((~g27472));
assign g13417 = ((~II20550));
assign g29132 = ((~II38139));
assign g28429 = (g17842&g28156);
assign g29140 = ((~II38163));
assign g23971 = (g18573&g23112);
assign g20109 = (g17878&g9504);
assign g24624 = ((~g23624)&(~g22555));
assign g11367 = ((~II18323));
assign g13412 = ((~II20535));
assign II17960 = ((~g6945));
assign g23140 = ((~g21825));
assign II32540 = ((~g24080))|((~II32538));
assign g4286 = ((~g2080));
assign g30203 = ((~g30027));
assign gbuf134 = (g1671);
assign g7782 = ((~g321));
assign II16880 = ((~g4203))|((~II16879));
assign II36138 = ((~g27547));
assign g15569 = ((~II21825));
assign II18282 = ((~g7923))|((~II18280));
assign II36230 = ((~g27583));
assign g29643 = ((~II39047));
assign gbuf25 = (g182);
assign g25210 = ((~g25000))|((~g3774));
assign g30482 = ((~g14067)&(~g30219));
assign g23395 = ((~g21973))|((~g22361));
assign g15324 = (g4609&g13196);
assign g30662 = ((~g16347)&(~g30469));
assign g13774 = ((~g12485));
assign g28375 = ((~II37280));
assign g20963 = ((~g19759)&(~g17715));
assign g20409 = ((~g17601));
assign II24444 = ((~g14148))|((~II24443));
assign g7335 = ((~g2827));
assign g30401 = ((~g29998)&(~g30128));
assign II31907 = ((~g23897));
assign g26577 = ((~g25436));
assign g28366 = ((~g15765)&(~g28116));
assign g3521 = ((~g1186));
assign g15671 = (g5242&g13273);
assign g5959 = ((~g876));
assign g13222 = ((~g9812));
assign g17664 = ((~II23748));
assign g28794 = ((~g28484)&(~g28009));
assign g10529 = (g5556&g5110);
assign g30767 = ((~II40555));
assign II35254 = ((~g26048));
assign g19821 = (g4705&g17776);
assign II14402 = ((~g1471));
assign II21505 = ((~g12952));
assign g20704 = ((~II27293));
assign g8330 = ((~II15532));
assign g29578 = ((~g28715)&(~g29188));
assign g16857 = ((~g15817)&(~g13023));
assign g26776 = ((~g26042)&(~g10024));
assign II36008 = ((~g26798));
assign g16189 = ((~g13043));
assign g24606 = ((~g24183)&(~g537));
assign II41135 = ((~g30975));
assign II31387 = ((~g22811));
assign g5162 = ((~g1294));
assign gbuf163 = (g1923);
assign II38833 = ((~g15962))|((~II38831));
assign g15432 = ((~II21694));
assign II26512 = ((~g16802));
assign g15003 = ((~g12269));
assign g5410 = ((~g3079));
assign g23271 = ((~II30266));
assign g5817 = (g1018&g1083);
assign II31733 = ((~g23603));
assign g29615 = (g29245&g11185);
assign g25948 = ((~g24564)&(~g24571));
assign II39863 = ((~g30278));
assign II20598 = ((~g13292));
assign g16105 = (g5622&g11797);
assign g23736 = ((~II30922));
assign g9365 = (g6314&g8056);
assign II21918 = ((~g11721));
assign g20769 = ((~II27358));
assign g24746 = (g15454&g24098);
assign g17924 = (g4930&g15547);
assign g8339 = (g6519&g903);
assign g20471 = ((~II26916));
assign g11983 = ((~g11284));
assign g12850 = ((~g8885));
assign g14684 = ((~II21262));
assign g22174 = ((~g19868)&(~g21593));
assign g22798 = (g18469&g21651);
assign II41132 = ((~g30974));
assign g29204 = ((~g15127)&(~g28915));
assign g23162 = ((~II29939));
assign g14592 = ((~g12263));
assign g30065 = ((~g29814)&(~g29817));
assign II23648 = ((~g15857));
assign g22809 = ((~g21850))|((~g21848))|((~g21879));
assign II38860 = ((~g29173));
assign g9639 = (g5438&g408);
assign II38125 = ((~g28425));
assign g30744 = (g30609&g20697);
assign g10213 = (g6751&g1255);
assign g20449 = ((~g17770));
assign g9187 = ((~g5803));
assign g24876 = (g24145&g20467);
assign II39053 = ((~g29546));
assign g15282 = (g4544&g13190);
assign g22047 = ((~g21313)&(~g19574));
assign g23136 = ((~g20878)&(~g10024));
assign g16371 = ((~g13095));
assign II35852 = ((~g26935));
assign g29162 = ((~II38229));
assign II24537 = ((~g14268))|((~g15118));
assign g29248 = (g28855&g8836);
assign g22627 = ((~II29223));
assign g22099 = ((~g21357)&(~g19651));
assign g23568 = ((~II30636));
assign II32170 = ((~g24231));
assign II29802 = ((~g21435));
assign g9173 = ((~II16465));
assign II18432 = ((~g6838));
assign g19725 = ((~II26154));
assign g7548 = ((~g2990));
assign g22421 = ((~g21012));
assign g16761 = ((~II22755));
assign II40703 = ((~g30649));
assign g23979 = ((~g23003)&(~g7009));
assign g26552 = ((~g25499));
assign g28674 = ((~II37569));
assign II38380 = ((~g28842))|((~II38378));
assign g22755 = ((~g21271)&(~g20842));
assign II15680 = ((~g7085));
assign g5826 = (g1718&g1749);
assign g28003 = ((~II36490));
assign g12747 = ((~g11421)&(~g8328)&(~g8385));
assign g27791 = ((~II36234));
assign II18464 = ((~g8620));
assign g19655 = (g4101&g17436);
assign g19454 = ((~g16611));
assign II18605 = ((~g9786));
assign II18438 = ((~g7265));
assign g9501 = ((~II16664));
assign g29074 = ((~II38035));
assign g9443 = ((~II16624));
assign II33570 = ((~g25065));
assign g25536 = ((~II33364));
assign g20900 = ((~g19648)&(~g17475));
assign g10846 = ((~g5799));
assign g23137 = ((~g17167)&(~g21218));
assign g17736 = (g4617&g15399);
assign II18160 = ((~g6783));
assign g26876 = ((~II35067));
assign II32642 = ((~g23348));
assign g13424 = ((~II20571));
assign g22997 = ((~g21706)&(~g21092));
assign g29901 = ((~g29687));
assign g25074 = ((~g24014))|((~g7303));
assign g15474 = ((~g12315));
assign II29259 = ((~g20925));
assign g25094 = ((~g23779));
assign g16878 = ((~II22855));
assign II35116 = ((~g26025));
assign g24613 = ((~g23592)&(~g22515));
assign g6134 = ((~II14647));
assign g7639 = ((~g3094));
assign g15499 = ((~II21758));
assign g10168 = (g3722&g4421);
assign II40904 = ((~g30733));
assign II14040 = ((~g2351));
assign g5249 = ((~g1961));
assign g13027 = ((~g9534))|((~g6912));
assign g7561 = ((~g1501));
assign g4913 = ((~g1063));
assign g19283 = (g14565)|(g16586);
assign g14131 = (g7727&g12961);
assign II36848 = ((~g27383));
assign II38838 = ((~g29357));
assign g29277 = ((~g28785));
assign g28149 = ((~g27667));
assign II33676 = ((~g24535));
assign g24358 = ((~II31748));
assign g5732 = ((~g1435));
assign II14755 = ((~g2821));
assign g16432 = (g2369&g12118);
assign g11874 = ((~g9808)&(~g9923)&(~g10059));
assign g30441 = (g30151&g11098);
assign g13902 = (g1928&g12829);
assign II37934 = ((~g28584));
assign g4520 = ((~g1395));
assign g10046 = (g3462&g1101);
assign II40991 = ((~g30794));
assign g20882 = ((~g19614)&(~g17408));
assign g5402 = ((~II13922));
assign g30133 = (g30067&g20799);
assign g18265 = ((~g14238));
assign g28978 = ((~g9150))|((~g28512));
assign g21284 = (g9356&g20269);
assign II19345 = ((~g10617));
assign II33586 = ((~g25052));
assign g7302 = ((~II14948));
assign II25778 = ((~g17145));
assign g8519 = (g6519&g876);
assign g23885 = ((~g22062));
assign g19629 = (g692&g18808);
assign g11812 = ((~II18990));
assign g30224 = (g30048&g9022);
assign g29634 = ((~II39020));
assign g28889 = ((~II37858));
assign g26739 = ((~II34824));
assign g11505 = ((~II18491));
assign II29280 = ((~g20936));
assign g26010 = ((~II33882));
assign II20535 = ((~g13359));
assign g24343 = ((~II31703));
assign g5985 = ((~g891));
assign g19740 = ((~II26171));
assign g3934 = ((~g176));
assign g29665 = ((~g29521)&(~g29289));
assign g27617 = ((~g27160));
assign g8494 = ((~II15696));
assign g29614 = (g29359&g11182);
assign g8387 = (g6232&g240);
assign II39423 = ((~g29666));
assign g12554 = ((~g8711));
assign g22717 = ((~II29405));
assign g28841 = (g27834&g28554);
assign g21610 = (g7522&g20490);
assign g4936 = ((~g1406));
assign g9580 = (g3410&g8209);
assign II40269 = ((~g30354));
assign g19087 = (g17215&g16540);
assign g28711 = (g10749&g28415);
assign II14280 = ((~g1491));
assign g28659 = (g27917&g13736);
assign g4251 = ((~g1115));
assign II29345 = ((~g20789));
assign g27428 = ((~II35768));
assign II35470 = ((~g26840));
assign II29421 = ((~g20983));
assign g14268 = ((~g12942));
assign g30824 = ((~II40724));
assign II23698 = ((~g15922));
assign g4780 = ((~g1263));
assign g30106 = (g29865&g11379);
assign g18404 = (g5343&g15794);
assign g22730 = ((~II29432));
assign g26659 = ((~g25334)&(~g17116));
assign g28849 = (g27850&g28616);
assign g19221 = (g18270)|(g18346);
assign g30388 = (g30229&g8918);
assign II31136 = ((~g22917));
assign g23075 = ((~g21628));
assign g11765 = ((~g10924));
assign g27073 = (g23381&g26634);
assign g28165 = ((~g27443));
assign g25118 = ((~II32844));
assign II30053 = ((~g22558));
assign g29572 = (g28802&g29397);
assign g18502 = ((~g14904));
assign g19043 = ((~II25192));
assign g19724 = (g2766&g18851);
assign g4982 = ((~g2208));
assign II36084 = ((~g27357));
assign II36256 = ((~g27527))|((~g15859));
assign II36708 = ((~g27324));
assign g26496 = ((~II34464));
assign g12070 = (g8018&g8766);
assign g16032 = (g12187&g10883);
assign g27872 = ((~II36337));
assign II29933 = ((~g22082));
assign g26858 = ((~II35017));
assign g25805 = ((~II33643));
assign g28033 = ((~II36560));
assign g20926 = ((~g19709)&(~g17599));
assign gbuf174 = (g2480);
assign II24521 = ((~g6435))|((~II24520));
assign g19849 = (g18014&g16126);
assign g30721 = ((~II40453));
assign g29178 = ((~g28848)&(~g28404));
assign g25658 = ((~II33482));
assign g27334 = ((~g27086)&(~g26449));
assign g22067 = ((~g21335)&(~g19605));
assign g22318 = ((~g20790));
assign II30155 = ((~g22737));
assign g22261 = ((~g20687));
assign g11321 = ((~II18271));
assign g10703 = ((~g3398))|((~g6678));
assign II37185 = ((~g27797));
assign II25802 = ((~g18265))|((~II25800));
assign II14742 = ((~g826));
assign g22518 = ((~II29064));
assign g10706 = ((~g3554))|((~g7162));
assign g13193 = ((~g9501));
assign II37050 = ((~g28081));
assign g21441 = ((~II27984));
assign g9724 = (g6574&g3972);
assign g3897 = ((~g2950));
assign g26713 = ((~II34746));
assign g15018 = ((~II21374));
assign g10208 = (g3410&g4504);
assign II32844 = ((~g23644));
assign g5115 = ((~g2651));
assign g22175 = (g16075)|(g20842);
assign g28066 = (g14596&g27555);
assign g21319 = (g9374&g20315);
assign II31577 = ((~g23782));
assign II24501 = ((~g6626))|((~II24500));
assign g26703 = ((~II34716));
assign g23560 = (g8206&g22428);
assign g21749 = (g3710&g20553);
assign g19818 = (g2052&g18902);
assign g15143 = (g4282&g13173);
assign II36912 = ((~g28024));
assign II39985 = ((~g30246));
assign g15510 = ((~II21769));
assign g22265 = (g21726&g12256);
assign II23341 = ((~g15784));
assign g17271 = ((~g16073)&(~g16106));
assign g30094 = (g29840&g11246);
assign g12960 = ((~g8997));
assign II35930 = ((~g26789));
assign II28825 = ((~g21882));
assign g21796 = ((~g19830)&(~g13004));
assign g22229 = (g21661&g12139);
assign g8504 = (g6369&g873);
assign g8183 = ((~g3188));
assign II26868 = ((~g17234));
assign g25250 = ((~g24822)&(~g23672));
assign g23559 = (g8203&g22425);
assign g21314 = (g9187&g20312);
assign II34153 = ((~g25234));
assign II32874 = ((~g24539));
assign g8088 = ((~g2549));
assign g28779 = ((~II37740));
assign g27292 = ((~g27026)&(~g26351));
assign II36150 = ((~g27569));
assign g30471 = ((~II40039));
assign g24745 = (g15454&g24096);
assign II35042 = ((~g26151))|((~g26145));
assign g11533 = ((~II18575));
assign g28440 = (g26092&g28162);
assign g13145 = ((~g9968))|((~g7488));
assign g17636 = (g4324&g16044);
assign g30325 = ((~II39818));
assign g24901 = (g24073&g18936);
assign g19762 = ((~II26195));
assign II33293 = ((~g25008));
assign g30023 = ((~g29548)&(~g29956));
assign g4475 = ((~g441));
assign II21520 = ((~g13067));
assign II33876 = ((~g25859));
assign II40481 = ((~g30676));
assign g18025 = ((~g14033));
assign g11831 = ((~g9648)&(~g9775)&(~g9904));
assign II23754 = ((~g16123));
assign g24430 = ((~g23393)&(~g10133));
assign g13429 = ((~II20586));
assign II35494 = ((~g26875));
assign g22249 = ((~g21699)&(~g20006));
assign g22341 = ((~g21169));
assign II14529 = ((~g3142));
assign g5918 = ((~g2379));
assign g30760 = (g30622&g22379);
assign g19634 = (g1326&g18810);
assign g24181 = ((~g16938)&(~g22220));
assign g14985 = ((~g11912));
assign g18743 = ((~g13648)&(~g11814));
assign II20553 = ((~g13290));
assign II38166 = ((~g29084));
assign g30097 = (g29849&g11271);
assign II28628 = ((~g21842));
assign II16453 = ((~g7936));
assign g12807 = ((~g8853));
assign II38936 = ((~g29212));
assign g20186 = (g13774&g13805&g13840&II26627);
assign g8551 = (g3566&g1573);
assign II17863 = ((~g7476));
assign g27732 = (g27492&g16758);
assign g18990 = (g13530&g16213);
assign II36105 = ((~g27517));
assign II23234 = ((~g9711))|((~II23233));
assign g21310 = (g9595&g20305);
assign II29724 = ((~g21851));
assign g20464 = ((~g17859));
assign g7958 = ((~g1175));
assign g22224 = (g21293&g16971);
assign II31895 = ((~g23846));
assign g30270 = ((~g16387)&(~g30104));
assign g21250 = ((~g19482)&(~g17183));
assign g28675 = ((~II37572));
assign g21557 = ((~II28087));
assign g18892 = ((~g15464));
assign g5810 = ((~g740));
assign g11151 = ((~II18067));
assign g23998 = ((~g22887))|((~g14044));
assign II21959 = ((~g13133));
assign g12154 = ((~g10383)&(~g10447)&(~g10511));
assign g19317 = (g16749&g3126);
assign g27432 = ((~II35772));
assign g13557 = ((~g12611))|((~g3410));
assign g30625 = ((~g30412)&(~g24660));
assign g24720 = ((~g23888)&(~g22759));
assign g27459 = ((~II35799));
assign II24178 = ((~g13873))|((~g9161));
assign g22906 = (g2924&g21927);
assign g23235 = ((~II30158));
assign g26732 = ((~II34803));
assign II21318 = ((~g12362));
assign II35301 = ((~g26037));
assign g17270 = ((~g16071)&(~g16104));
assign g26636 = ((~g25767));
assign II32854 = ((~g24092));
assign g23997 = ((~g22887))|((~g14048));
assign g21799 = (g16505)|(g20538)|(g18994)|(II28318);
assign g10235 = ((~II17209));
assign g25619 = (g14497&g25111);
assign g29935 = ((~II39407));
assign g10077 = (g7085&g4298);
assign g23455 = ((~II30489));
assign g12926 = (g9676)|(g3554);
assign g20246 = (g16778&g16974&g16743);
assign II39782 = ((~g30054));
assign g18691 = ((~g14885));
assign g19558 = (g8056&g17252);
assign g19148 = (g17202&g16817);
assign g21063 = ((~g19913)&(~g15710));
assign g20611 = ((~II27158));
assign g5932 = ((~g813));
assign g26362 = (g4891&g25640);
assign g25122 = ((~II32854));
assign g21792 = ((~g20255))|((~g7085));
assign g10407 = (g5556&g2513);
assign g13865 = (g548&g12748);
assign g24373 = ((~II31793));
assign g20281 = ((~g17243));
assign II35124 = ((~g26107))|((~II35123));
assign g22962 = ((~g21763));
assign g15774 = ((~II22022));
assign II30860 = ((~g22106));
assign II21407 = ((~g13039));
assign g16350 = (g981&g11985);
assign g24854 = ((~II32499))|((~II32500));
assign II40131 = ((~g30493));
assign II29697 = ((~g21082));
assign II18226 = ((~g5668));
assign g11749 = ((~II18929));
assign II20347 = ((~g10787));
assign g13186 = ((~g9446));
assign g29679 = ((~g29549)&(~g29329));
assign g7876 = ((~II15191))|((~II15192));
assign g16894 = (g7156&g14959);
assign g28101 = ((~II36738));
assign g24941 = ((~g23526));
assign II32153 = ((~g24223));
assign g12307 = (g7919&g8853);
assign g4962 = ((~g1970));
assign g24663 = ((~g24183)&(~g532));
assign g12048 = ((~g10219)&(~g10304)&(~g10381));
assign g24711 = ((~g24183)&(~g536));
assign II16044 = ((~g5397));
assign II31919 = ((~g23524));
assign g5876 = ((~g2180));
assign II37038 = ((~g28038));
assign II36240 = ((~g27603));
assign g22655 = ((~II29271));
assign g7872 = ((~g2874));
assign g19840 = (g679&g18910);
assign g21952 = ((~II28482));
assign g9026 = (g5438&g7610);
assign g29050 = ((~II38007));
assign g10095 = ((~II17060))|((~II17061));
assign g29241 = (g9711&g28823);
assign g23670 = ((~II30816));
assign II37083 = ((~g28102));
assign II30925 = ((~g22127));
assign g22692 = ((~II29348));
assign II25750 = ((~g2129))|((~g18390));
assign g29345 = ((~g28339)&(~g28726));
assign II27672 = ((~g20545));
assign g16993 = (g7576&g15322);
assign g27785 = ((~II36224));
assign II25474 = ((~g18885));
assign II24530 = ((~g6707))|((~g14355));
assign g30155 = ((~g30015));
assign g23055 = ((~II29802));
assign g17936 = (g4942&g15557);
assign g11444 = ((~II18408));
assign II40294 = ((~g30470));
assign g25554 = ((~II33382));
assign g22289 = (g780&g21565);
assign II32569 = ((~g24082))|((~II32567));
assign II15222 = ((~g3151));
assign II35521 = ((~g26883));
assign g26674 = (g25291&g21090);
assign g17463 = (g4150&g15136);
assign g5893 = ((~g125));
assign g25220 = ((~g24762)&(~g23573));
assign II39797 = ((~g30307));
assign g19153 = ((~g17381)&(~g15093));
assign II38378 = ((~g28845))|((~g28842));
assign g13070 = ((~II20117));
assign g17132 = ((~g15981)&(~g15971)&(~g15952));
assign II23821 = ((~g14337));
assign II26940 = ((~g17383));
assign g27736 = ((~g27396)&(~g26962));
assign g20793 = ((~II27382));
assign g8707 = ((~II15909));
assign g27956 = ((~II36423));
assign g24569 = (g767&g23455);
assign II39776 = ((~g30066));
assign g8879 = ((~II16147));
assign II28564 = ((~g21385));
assign g18195 = ((~II24195))|((~II24196));
assign g13941 = (g7635&g12859);
assign g4828 = ((~g1822));
assign g26616 = ((~g13860)&(~g25310));
assign g20632 = ((~II27221));
assign g16493 = ((~II22581));
assign II25829 = ((~g2138))|((~g18314));
assign g29101 = ((~II38094));
assign II31676 = ((~g23517));
assign g30035 = ((~II39540))|((~II39541));
assign g20827 = ((~II27416));
assign g21129 = (g20273&g12302);
assign g25286 = (g24668&g8752);
assign g9912 = (g5473&g4144);
assign g27134 = ((~g26175));
assign g8813 = ((~II16027));
assign g30511 = ((~II40113));
assign II25921 = ((~g2151))|((~g18526));
assign g8266 = ((~II15466));
assign II22512 = ((~g13635));
assign g23621 = ((~II30741));
assign g16840 = ((~g15878));
assign II27107 = ((~g19249));
assign g28582 = ((~g27820));
assign g29553 = (g29223&g29386);
assign II39168 = ((~g29623));
assign g25865 = ((~II33711));
assign g29680 = ((~g29553)&(~g29330));
assign II35961 = ((~g26825));
assign g26953 = ((~II35136));
assign II34791 = ((~g26489));
assign g22480 = ((~II29026));
assign g29100 = ((~II38091));
assign g13232 = ((~g9895));
assign g11905 = ((~g9920)&(~g10056)&(~g10144));
assign g21044 = ((~g19885)&(~g18059));
assign g16201 = ((~g13073));
assign g28058 = (g27604&g10052);
assign g10218 = (g7162&g4520);
assign g25634 = ((~II33457));
assign g12942 = ((~g8507)&(~g8522)&(~g8537));
assign g15244 = (g7852&g12695);
assign g23317 = ((~II30404));
assign g27568 = (g24004&g27172);
assign g30555 = ((~II40245));
assign g21523 = (g15296&g20465);
assign g13386 = ((~II20483));
assign II29672 = ((~g21074));
assign II38878 = ((~g29185));
assign g23079 = ((~g21640));
assign g21926 = (g19354&g13011);
assign g562 = ((~II13089));
assign g22941 = ((~g8305))|((~g21751));
assign g25343 = ((~g24975)&(~g5623));
assign g9898 = ((~II16900));
assign g22748 = ((~II29478));
assign II16873 = ((~g6102));
assign II28090 = ((~g20008));
assign II35689 = ((~g26878));
assign g21167 = ((~g20159)&(~g20189));
assign g29916 = ((~g24712)&(~g29726));
assign II36894 = ((~g28022));
assign g8840 = ((~II16074));
assign g13870 = (g7582&g12768);
assign II40970 = ((~g30782));
assign g7967 = ((~g2966));
assign g12332 = ((~g10829));
assign g21095 = ((~g20012)&(~g20049)&(~g20084));
assign g25646 = ((~II33469));
assign g30708 = ((~g14212)&(~g30396));
assign g13212 = ((~g9734));
assign g10477 = (g7426&g5015);
assign g22338 = ((~g20806));
assign g23905 = ((~g22046));
assign II40078 = ((~g30263));
assign g19225 = (g18383)|(g18561);
assign II17698 = ((~g6711));
assign g24695 = (g13576&g24134);
assign g13673 = ((~II20886));
assign g11894 = ((~g11141));
assign g30306 = ((~II39761));
assign g23501 = ((~II30547));
assign g27724 = ((~g27254)&(~g10340));
assign g12768 = ((~g8829));
assign II38602 = ((~g29016));
assign II20625 = ((~g13367));
assign II30122 = ((~g22827));
assign II32607 = ((~g18038))|((~g24090));
assign II36604 = ((~g27296));
assign II16082 = ((~g5401));
assign g11868 = ((~g11098));
assign II31460 = ((~g23728));
assign g29209 = ((~g15196)&(~g28936));
assign II28034 = ((~g19173));
assign g7579 = ((~g1877));
assign g11779 = ((~g10906));
assign g20922 = ((~g19698)&(~g17577));
assign II29174 = ((~g20899));
assign II19432 = ((~g10653));
assign II27206 = ((~g20471));
assign g10127 = ((~II17103));
assign g12105 = ((~g11456));
assign g27011 = ((~g24916)&(~g26026));
assign g15476 = (g4929&g13221);
assign g10293 = (g6678&g4626);
assign g22477 = ((~II29023));
assign g23680 = (g4307&g22570);
assign g26513 = ((~g25389))|((~g2133));
assign g26433 = ((~II34392));
assign II24485 = ((~g14541))|((~g9391));
assign g13173 = ((~g9338));
assign g23598 = (g4038&g22484);
assign g18666 = (g14849&g13687&g13714&g16302);
assign g5092 = ((~g2098));
assign g11771 = (g554&g8622);
assign g30735 = (g30629&g22268);
assign II18749 = ((~g8779));
assign II28305 = (g20197)|(g20177)|(g20145);
assign g27327 = ((~g27077)&(~g26432));
assign II34476 = ((~g25201));
assign g22953 = ((~g20700)&(~g7595));
assign g26272 = ((~g25973)&(~g16423));
assign g16136 = (g5640&g11819);
assign g15834 = ((~g12611))|((~g6369));
assign g8822 = ((~g4602));
assign g20355 = ((~g17422));
assign II27361 = ((~g19390));
assign g29799 = ((~II39249));
assign g25566 = (g24843)|(g23143);
assign g26799 = ((~g26158)&(~g25453));
assign g28356 = ((~g15680)&(~g28086));
assign g28229 = ((~II36936));
assign g5352 = ((~g737));
assign g13068 = ((~g9968))|((~g7488));
assign II35944 = ((~g27078))|((~g14904));
assign g18861 = ((~g15363));
assign g23662 = ((~II30800));
assign g4130 = ((~g846));
assign g25540 = ((~II33368));
assign g21711 = ((~g19830)&(~g15780));
assign g23099 = ((~g21180)&(~g21208));
assign g28456 = (g28141&g9351);
assign g16342 = (g5894&g11968);
assign g28647 = ((~g27959));
assign II22533 = ((~g14795));
assign II13095 = ((~g1943));
assign II31520 = ((~g23683));
assign g29534 = (g29206&g29374);
assign g8321 = ((~II15523));
assign g27216 = ((~II35485));
assign II35503 = ((~g26896));
assign II26078 = ((~g16835));
assign g5657 = ((~II14113));
assign II24037 = ((~g14016))|((~II24036));
assign g27448 = (g2766&g27142);
assign g6163 = ((~g1365));
assign II18052 = ((~g6232));
assign g17381 = (g8250&g16001);
assign g10615 = (g3522&g5243);
assign g11354 = ((~II18308));
assign g30355 = (g30207&g8421);
assign g17913 = ((~II23959))|((~II23960));
assign II36574 = ((~g27289));
assign II25141 = ((~g18970));
assign g11432 = ((~II18396));
assign g27042 = (g21996&g26608);
assign g13637 = ((~g11703));
assign g19121 = ((~g16682))|((~g16697));
assign g19703 = (g4240&g17517);
assign g10826 = ((~II17673));
assign g13310 = ((~g11481)&(~g11332)&(~g11190)&(~g11069));
assign II19921 = ((~g8563));
assign g24867 = (g666&g23779);
assign g20746 = ((~II27335));
assign g27146 = ((~g26358));
assign II14073 = ((~g2574));
assign g28083 = ((~II36690));
assign g23839 = ((~II31077));
assign II25847 = ((~g771))|((~II25846));
assign g26289 = (g4595&g25527);
assign g25039 = ((~g23803))|((~g7265));
assign II31065 = ((~g22166));
assign g29549 = (g26043&g29384);
assign g19000 = ((~II25084));
assign g28155 = ((~g27404));
assign g11724 = ((~g9822))|((~g3678));
assign g26341 = ((~II34296));
assign g10016 = ((~II16984));
assign g27358 = (g749&g26846);
assign g13279 = ((~g10161));
assign g26956 = ((~II35141));
assign g22296 = ((~g20754));
assign g13309 = ((~g10276));
assign g20435 = ((~g17701));
assign g6782 = ((~II14831));
assign g9401 = ((~II16598));
assign g28854 = (g27892&g28629);
assign II26654 = (g14936&g18815&g13774);
assign g12912 = ((~g8484)&(~g8500)&(~g8515));
assign g4375 = ((~g1110));
assign g16457 = (g5831&g13391);
assign g23202 = ((~II30059));
assign g12159 = ((~g8354));
assign II40733 = ((~g30659));
assign g29062 = ((~g9310))|((~g28540));
assign II38689 = ((~g29325));
assign g29366 = ((~g28906));
assign g13043 = ((~g10789));
assign g8472 = (g3566&g1609);
assign g18124 = ((~g14551)&(~g16058));
assign II27827 = ((~g19896));
assign II37784 = ((~g28567));
assign II40835 = ((~g30816));
assign II21647 = ((~g11695));
assign g10220 = (g6980&g4526);
assign g24129 = ((~g22477));
assign II35695 = ((~g26887));
assign g29272 = ((~g28768));
assign g27585 = ((~g26950)&(~g24739));
assign g24453 = ((~g23694))|((~g3462));
assign g9446 = ((~II16627));
assign g12418 = ((~g10729)&(~g10748)&(~g10764));
assign II30976 = ((~g22142));
assign II14877 = ((~g1309));
assign g30260 = ((~g16322)&(~g30094));
assign II25303 = ((~g17151));
assign II27113 = ((~g19689));
assign g9094 = (g6713&g7679);
assign g16728 = ((~g14910));
assign g22770 = (g14414&g21628);
assign II25030 = ((~g8029))|((~g13507));
assign g21699 = (g3710&g20518);
assign II14014 = ((~g499));
assign g23689 = (g6513&g23001);
assign II37593 = ((~g28443));
assign g18878 = ((~g15429));
assign g8179 = ((~g3062));
assign g13105 = ((~g9822))|((~g7230));
assign g30861 = ((~II40835));
assign g30312 = ((~II39779));
assign II19654 = ((~g10805));
assign g11547 = ((~II18617));
assign g16954 = ((~g13589));
assign g20118 = (g13687&g13714&g13791&II26564);
assign II18680 = ((~g8973));
assign g24126 = ((~g20928))|((~g22199));
assign g23741 = (g22708&g17667);
assign g18038 = ((~II24071));
assign g24464 = ((~g23955))|((~g3494));
assign g28387 = (g1426&g27787);
assign g30703 = ((~g14022)&(~g30391));
assign gbuf98 = (g1012);
assign II30701 = ((~g22057));
assign II27324 = ((~g19358));
assign g20105 = ((~II26545));
assign g30000 = (g10767&g29930);
assign g23045 = ((~g21577));
assign g5897 = ((~g267));
assign g12050 = ((~g10222)&(~g10309)&(~g10387));
assign g11066 = ((~II17984));
assign g12275 = ((~g8303));
assign II25810 = ((~g767))|((~II25809));
assign g11897 = ((~g9907)&(~g10043)&(~g10118));
assign g19531 = (g16884&g16722&g14776);
assign g18943 = ((~g15655));
assign g21461 = ((~g19957));
assign g27287 = ((~g27021)&(~g26342));
assign g16853 = ((~g15801)&(~g13009));
assign g16041 = ((~g12762));
assign g13465 = ((~II20694));
assign g10436 = (g6912&g4902);
assign II16900 = ((~g6486));
assign II26464 = (g18370&g18296&g18206);
assign g30015 = ((~g29527)&(~g29948));
assign II35437 = ((~g27183));
assign II24655 = ((~g6190))|((~g14592));
assign II27772 = (g19314&g19501&g19480);
assign g26189 = ((~g25952));
assign g8847 = ((~II16089));
assign g23936 = ((~g22812))|((~g13922));
assign g24301 = ((~II31577));
assign II32577 = ((~g24089))|((~II32575));
assign II30083 = ((~g22676));
assign II14984 = ((~g2625));
assign g15437 = (g4869&g13214);
assign II24513 = ((~g13992))|((~II24512));
assign g27410 = ((~II35750));
assign g22743 = ((~II29465));
assign g26584 = ((~g25590));
assign g24101 = ((~g22415));
assign gbuf14 = (g2842);
assign II24381 = ((~g6212))|((~II24380));
assign g12057 = ((~g10228)&(~g10313)&(~g10391));
assign II30074 = ((~g22648));
assign g19511 = ((~g16788));
assign g26921 = ((~II35116));
assign g25438 = ((~g24982));
assign II25633 = ((~g65))|((~g17640));
assign g26599 = ((~g25637));
assign g24593 = ((~II32167));
assign g8993 = ((~II16309));
assign g29413 = ((~II38620));
assign g23262 = ((~II30239));
assign II40814 = ((~g30731));
assign II39151 = ((~g29617));
assign g12447 = ((~II19615));
assign g15486 = (g4797&g12822);
assign g15376 = ((~II21638));
assign g22702 = ((~II29366));
assign g8910 = ((~II16196));
assign g21048 = ((~g19889)&(~g18062));
assign g19180 = ((~II25395));
assign II22626 = ((~g15151));
assign g29694 = ((~II39136));
assign g29375 = ((~g28955));
assign g15931 = ((~g12711))|((~g6838));
assign g10419 = ((~II17373));
assign II32184 = ((~g23497));
assign II16074 = ((~g5399));
assign g18275 = ((~g14171));
assign II24388 = ((~g6421))|((~II24387));
assign II38635 = ((~g29305));
assign g11841 = ((~g11048));
assign g28345 = ((~g15527)&(~g28028));
assign g8632 = ((~II15822));
assign g30800 = ((~II40654));
assign g9138 = (g5556&g7806);
assign II39017 = ((~g29542));
assign II23448 = ((~g15834));
assign g11166 = ((~II18082));
assign g23204 = ((~II30065));
assign g13894 = ((~g11806));
assign g26911 = ((~g25569))|((~g26283));
assign II30179 = ((~g22657));
assign g20383 = ((~g17503));
assign g17360 = ((~II23448));
assign g17450 = (g4124&g15115);
assign II14799 = ((~g551));
assign II37041 = ((~g28060));
assign II23463 = ((~g15812));
assign g24793 = (g9857&g24144);
assign g8259 = ((~II15445));
assign g21292 = (g9453&g20281);
assign g18882 = ((~g15449));
assign g23070 = ((~g21140)&(~g21173));
assign g12064 = ((~g11398));
assign g12150 = ((~g8341));
assign g13624 = ((~II20852));
assign II20873 = ((~g12482));
assign g15992 = ((~g12886))|((~g6678));
assign g28963 = ((~g28664)&(~g13365));
assign II20697 = ((~g13369));
assign g22846 = ((~g8278))|((~g21660));
assign g27056 = (g22069&g26622);
assign g28758 = ((~g15126)&(~g28451));
assign II34198 = ((~g25245));
assign g17830 = ((~II23894))|((~II23895));
assign g29094 = ((~II38077));
assign g12969 = ((~g9010));
assign g10074 = (g7230&g4289);
assign II38011 = ((~g28584));
assign II15899 = ((~g5626));
assign g29418 = ((~II38635));
assign g19478 = ((~II25914))|((~II25915));
assign g5646 = ((~g213));
assign g3987 = ((~g2224));
assign g25772 = ((~g24624)&(~g24520));
assign II33154 = ((~g25005));
assign g19754 = (g2026&g18861);
assign g18324 = ((~g14329));
assign g19882 = (g18131&g16177);
assign II25108 = ((~g18969));
assign g18871 = ((~g15396));
assign II39532 = ((~g29915))|((~g29917));
assign g9082 = (g3650&g1870);
assign g21378 = (g9507&g20378);
assign II32634 = ((~g18131))|((~II32633));
assign g26114 = ((~II34009));
assign g8391 = ((~II15593));
assign g23209 = ((~II30080));
assign g15573 = (g4976&g12863);
assign g24810 = (g9857&g24160);
assign II37982 = ((~g28501));
assign g19671 = (g4159&g17468);
assign g16285 = (g2590&g11921);
assign II18031 = ((~g7195));
assign g13669 = ((~g13229));
assign II30296 = ((~g22723));
assign g9484 = ((~II16653));
assign II33732 = ((~g24473));
assign g23583 = (g3978&g22467);
assign g27149 = ((~g23462)&(~g26060));
assign g27163 = ((~II35364));
assign II38046 = ((~g28348));
assign g28447 = ((~II37400));
assign g26642 = ((~g25793));
assign g24235 = ((~g17062)&(~g22305));
assign g14736 = ((~g11957));
assign g27371 = (g2129&g26861);
assign g17330 = ((~II23418));
assign II22962 = ((~g9161))|((~g13885));
assign g26983 = ((~II35172));
assign II18728 = ((~g8878));
assign g24213 = ((~g16988)&(~g22245));
assign g30697 = (g30383&g11011);
assign g5901 = ((~g939));
assign g12302 = ((~II19472));
assign g21235 = ((~g19281)&(~g19269));
assign g30561 = ((~II40263));
assign g14584 = ((~g11811));
assign g5710 = (g331&g381);
assign II30314 = ((~g22772));
assign g5871 = ((~g1685));
assign g28763 = ((~g15160)&(~g28456));
assign g28724 = (g28551&g16725);
assign g24382 = ((~II31820));
assign g11968 = ((~g11265));
assign g6944 = ((~II14865));
assign g25335 = ((~g24832));
assign g19165 = ((~g17526)&(~g15264));
assign g6290 = ((~g1332));
assign g24723 = (g13605&g24168);
assign g29009 = ((~g28669)&(~g28320));
assign g24774 = (g2052&g24127);
assign g14086 = ((~g11938));
assign g24336 = ((~II31682));
assign g29358 = ((~g29120));
assign g18834 = ((~g15240));
assign g28061 = ((~II36630));
assign g5556 = ((~II14040));
assign II37191 = ((~g27792));
assign g5764 = ((~g918));
assign g12210 = ((~g8400));
assign g10196 = (g3306&g435);
assign g22169 = ((~g21448)&(~g19782));
assign II35868 = ((~g26812));
assign g20633 = ((~g20164))|((~g3254));
assign g13141 = ((~g9146));
assign g19100 = (g17220&g16596);
assign g18765 = ((~g14991));
assign g7623 = ((~g314));
assign II32724 = ((~g23913))|((~g14514));
assign g25868 = ((~II33714));
assign g24109 = ((~g20904))|((~g22190));
assign g20596 = ((~II27113));
assign g10171 = (g3722&g4430);
assign g5920 = (g2406&g2471);
assign II29575 = ((~g21042));
assign g28252 = ((~II37005));
assign g30217 = (g30036&g8955);
assign g27553 = ((~II35953));
assign II23567 = ((~g15839));
assign g27534 = (g23974&g27155);
assign g23798 = (g7079&g23031);
assign II18701 = ((~g11471));
assign g19150 = (g17189&g8602);
assign II40667 = ((~g30637));
assign II40320 = ((~g30341));
assign g23082 = ((~g21647));
assign g20607 = ((~II27146));
assign g18587 = ((~II24684));
assign II15958 = ((~g3878));
assign II23968 = ((~g9248))|((~II23966));
assign g24514 = ((~g23798)&(~g22682));
assign II35772 = ((~g26772));
assign g6098 = ((~II14609));
assign g23187 = ((~II30014));
assign g12263 = ((~g10524)&(~g10586)&(~g10627));
assign g30163 = ((~g30017));
assign II30568 = ((~g23114));
assign II19485 = ((~g10617));
assign II29975 = ((~g22641));
assign g23186 = ((~II30011));
assign g29786 = ((~g29486)&(~g29239));
assign II25129 = ((~g16813));
assign g12487 = ((~g10108)&(~g10198)&(~g10283));
assign g28008 = (g27590&g9770);
assign g26434 = ((~II34395));
assign II15978 = ((~g7303));
assign II40179 = ((~g30498));
assign g22831 = ((~g21285)&(~g20858));
assign g26885 = ((~g26140)&(~g22319));
assign g21660 = ((~II28190))|((~II28191));
assign II26596 = (g18708&g18735&g18765);
assign g20314 = ((~g13646)&(~g16855));
assign g17599 = (g4383&g15268);
assign g19174 = ((~II25383));
assign II21286 = ((~g11678));
assign g24817 = ((~II32392))|((~II32393));
assign g25338 = ((~g24860));
assign g13130 = ((~g9140));
assign g27824 = ((~g6087)&(~g27632)&(~g25399));
assign II35919 = ((~g26938));
assign g29877 = ((~g29681));
assign II28229 = ((~g20067));
assign II24394 = ((~g15995));
assign II24626 = ((~g14252))|((~II24624));
assign II23074 = ((~g9293))|((~g13856));
assign g4651 = ((~g1128));
assign II28051 = ((~g20025));
assign g28094 = (g27617&g10179);
assign gbuf201 = (g2597);
assign II25732 = ((~g758))|((~II25731));
assign II27212 = ((~g20498));
assign g8221 = ((~g860));
assign g10476 = (g7488&g5012);
assign g26532 = ((~g25979)&(~g17100));
assign g9383 = (g6369&g8068);
assign II38695 = ((~g29326));
assign g20468 = ((~g17871));
assign g10444 = (g3494&g1279);
assign g6027 = ((~g2339));
assign g21016 = ((~g19847)&(~g17925));
assign g18989 = ((~II25057));
assign g30070 = ((~g29827)&(~g29833));
assign g26600 = ((~g25640));
assign g20612 = ((~II27161));
assign g4641 = ((~g1033));
assign g10804 = ((~II17649));
assign g18606 = ((~II24710))|((~II24711));
assign g20459 = ((~II26898));
assign II40889 = ((~g30825));
assign g20903 = ((~g19662)&(~g17510));
assign g21021 = ((~g19853)&(~g17949));
assign g22217 = ((~g21928));
assign g28105 = (g27613&g10235);
assign II24913 = ((~g15800));
assign g9759 = (g3254&g4000);
assign II17966 = ((~g7015));
assign g19060 = ((~II25243));
assign gbuf91 = (g1054);
assign II17872 = ((~g7539));
assign gbuf52 = (g551);
assign g21959 = ((~II28503));
assign g11376 = ((~II18332));
assign II22828 = ((~g14514));
assign g30921 = (g10773&g30791);
assign g10371 = (g6912&g4766);
assign g5409 = ((~II13943));
assign II31628 = ((~g23621));
assign g19921 = ((~g16639))|((~g9928));
assign II24194 = ((~g13927))|((~g15188));
assign g20640 = (g4809&g19064);
assign II16150 = ((~g3900));
assign g22074 = ((~g21338)&(~g19617));
assign g8440 = ((~II15642));
assign g27047 = (g23344&g26613);
assign g28783 = ((~g28466)&(~g27968));
assign g20148 = (g13724&g13764&g13819&II26596);
assign II25721 = ((~g74))|((~g18341));
assign g4544 = ((~g1804));
assign II31688 = ((~g24035));
assign g20875 = ((~g19584)&(~g17352));
assign g4647 = ((~g1071));
assign II39622 = ((~g30052));
assign g17506 = (g6675&g16023);
assign g27667 = ((~II36046));
assign II33867 = ((~g25833));
assign g9462 = (g6519&g8141);
assign g21995 = ((~II28550));
assign g6180 = ((~g692));
assign g17222 = ((~g15998)&(~g16003));
assign g27718 = ((~g27251)&(~g10133));
assign g28321 = ((~g27742)&(~g10133));
assign g16616 = ((~II22663));
assign g21270 = (g20357&g15080);
assign II31601 = ((~g23562));
assign g14718 = ((~II21277));
assign g10465 = (g7230&g4979);
assign g23605 = (g4067&g22497);
assign II30552 = ((~g23097));
assign g21361 = (g9150&g20362);
assign II39404 = ((~g29661));
assign g8554 = (g3566&g1654);
assign g19334 = ((~II25722))|((~II25723));
assign g8545 = (g6838&g2342);
assign g8098 = ((~g3051));
assign g23633 = ((~II30763));
assign g24418 = ((~II31928));
assign g9248 = ((~g5859));
assign g9479 = (g6783&g8150);
assign g22824 = ((~II29603));
assign g26663 = (g25274&g21066);
assign g5543 = ((~g3087));
assign II37725 = ((~g28540));
assign II36676 = ((~g27315));
assign II32102 = ((~g24182));
assign g28391 = ((~II37323))|((~II37324));
assign g9756 = ((~g5504));
assign g15820 = ((~g12565))|((~g6232));
assign gbuf208 = (g2549);
assign g10461 = (g7358&g4967);
assign g5255 = ((~g1988));
assign II23451 = ((~g13497));
assign g24826 = (g12974&g24167);
assign g8835 = ((~II16065));
assign g14366 = ((~g12090));
assign gbuf177 = (g2529);
assign g22640 = ((~II29246));
assign g27120 = ((~g26560)&(~g17001));
assign g11991 = ((~g10146)&(~g10218)&(~g10303));
assign g10118 = (g3410&g4366);
assign g17543 = (g4289&g15228);
assign II34659 = ((~g26190));
assign II24076 = ((~g14414))|((~g9277));
assign II19702 = ((~g10125));
assign II36738 = ((~g27331));
assign g22202 = (g21626&g21036);
assign g17057 = ((~g13519));
assign g30928 = ((~II41024));
assign g30540 = ((~II40200));
assign g27230 = ((~II35527));
assign g25133 = ((~II32877));
assign g30267 = ((~g16380)&(~g30101));
assign g28709 = (g28400&g22261);
assign g22623 = ((~II29215));
assign II38641 = ((~g29249));
assign II31904 = ((~g23873));
assign II33421 = ((~g25043));
assign g21842 = ((~g13609)&(~g19150));
assign g25368 = ((~g24778));
assign II37324 = ((~g27855))|((~II37322));
assign g17903 = ((~II23954));
assign g21457 = ((~II28000));
assign g22789 = ((~g21278)&(~g20850));
assign g30470 = ((~g14023)&(~g30218));
assign II23958 = ((~g6513))|((~g14171));
assign g10048 = (g6713&g4251);
assign g30656 = ((~g16310)&(~g30460));
assign g22408 = ((~g20986));
assign g22367 = ((~g21242));
assign g30079 = (g29823&g10988);
assign g28540 = (g26497)|(g27743);
assign II37176 = ((~g27927));
assign g25402 = ((~II33232));
assign g29156 = ((~II38211));
assign II31589 = ((~g23856));
assign g19041 = ((~II25186));
assign g21700 = ((~II28229));
assign g16515 = ((~g14244));
assign II40071 = ((~g30261));
assign g24962 = ((~g23764));
assign g13449 = ((~II20646));
assign g27768 = ((~g27568)&(~g27110));
assign g30456 = ((~II40016));
assign g17887 = ((~II23942))|((~II23943));
assign g28398 = (g7769&g27817);
assign g13882 = ((~g11790));
assign g18863 = ((~g15379));
assign g17601 = ((~II23689));
assign II38975 = ((~g29348));
assign II28133 = (g18025&g18453&g18110);
assign g20127 = ((~g18623));
assign g30126 = ((~II39641));
assign g5272 = ((~g2657));
assign g24110 = ((~g22437));
assign g11465 = ((~II18429));
assign g12231 = ((~g10473)&(~g10532)&(~g10591));
assign g4098 = ((~g156));
assign g22034 = ((~g21302)&(~g19561));
assign g22240 = ((~g20652));
assign g23866 = (g22971&g9819);
assign II35890 = ((~g26815));
assign g22015 = (g1672&g21217);
assign g28431 = (g26092&g28158);
assign g21786 = ((~g14577))|((~g15441))|((~g19942))|((~g19931));
assign g18962 = ((~g15731));
assign II20959 = ((~g11713));
assign g27095 = (g5173&g26442);
assign g30299 = ((~g13499)&(~g29996));
assign g30570 = ((~g30404));
assign g19113 = ((~II25308));
assign g9505 = ((~g6227));
assign g19480 = ((~II25922))|((~II25923));
assign g26542 = ((~g25472));
assign g18877 = ((~g15426));
assign II40170 = ((~g30483));
assign g10995 = ((~II17898));
assign II23105 = ((~g14052))|((~II23103));
assign g6887 = ((~g2584));
assign II17978 = ((~g7795));
assign g11863 = ((~g9774)&(~g9902)&(~g10035));
assign g26191 = ((~II34099));
assign II23253 = ((~g13741));
assign g5998 = ((~g2336));
assign g13858 = ((~g11603));
assign II22974 = ((~g13962))|((~II22972));
assign II14811 = ((~g623));
assign II13907 = ((~g1030));
assign II17677 = ((~g6517));
assign II39899 = ((~g30288));
assign g21778 = ((~g19494)&(~g18121)&(~g14309));
assign g7970 = ((~II15277))|((~II15278));
assign g21393 = (g9264&g20389);
assign g29525 = (g29195&g29366);
assign g10595 = (g7391&g2673);
assign II21769 = ((~g11705));
assign g25030 = ((~g23923))|((~g6643));
assign g30468 = ((~g14007)&(~g30217));
assign g22886 = ((~g16164)&(~g20858)&(~g21285));
assign g29648 = ((~II39062));
assign gbuf159 = (g1855);
assign II18399 = ((~g6519));
assign g25838 = ((~II33680));
assign g8894 = ((~II16166));
assign II36673 = ((~g27314));
assign g12076 = ((~g11414));
assign II15964 = ((~g7554));
assign II22768 = ((~g14691));
assign g6638 = ((~g3103));
assign g5978 = ((~II14446));
assign g24066 = ((~II31286));
assign g15336 = (g4492&g12752);
assign g20555 = ((~II26990));
assign II29087 = ((~g20728));
assign g19214 = (g18383)|(g18458);
assign g23304 = ((~II30365));
assign g29453 = ((~II38740));
assign II16292 = ((~g5426));
assign g15524 = ((~g12333));
assign g20013 = (g17720&g12848);
assign g18831 = ((~g15228));
assign g19813 = (g4677&g17758);
assign g30538 = ((~II40194));
assign g27254 = ((~g26968)&(~g26231));
assign g15801 = (g7856&g13351);
assign g30515 = ((~II40125));
assign II13919 = ((~g1045));
assign II39843 = ((~g30273));
assign g23192 = ((~II30029));
assign II34204 = ((~g25247));
assign g11816 = (g7869&g8655);
assign g20979 = ((~g19786)&(~g17775));
assign g19385 = (g16954&g16619&g14423);
assign g12995 = ((~g8545)&(~g8558)&(~g8567));
assign II17666 = ((~g6430));
assign g6642 = ((~II14799));
assign II29957 = ((~g22585));
assign II30838 = ((~g22100));
assign g23193 = ((~II30032));
assign II36300 = ((~g27382))|((~g27379));
assign g22304 = ((~g20766));
assign g12923 = ((~g10147)&(~g6421));
assign g21473 = ((~II28009));
assign g22021 = ((~g21609))|((~g21634));
assign g13158 = ((~g9242));
assign g10184 = (g7488&g4447);
assign g13242 = ((~g9962));
assign g19755 = (g4421&g17621);
assign g22734 = ((~II29442));
assign g24349 = ((~II31721));
assign g26216 = ((~II34146));
assign g25880 = ((~II33726));
assign g16692 = ((~g14752)&(~g12514));
assign g18312 = ((~g14554));
assign g29312 = (g29049&g28955);
assign g22763 = ((~II29509));
assign g28339 = (g28059&g19498);
assign g11976 = ((~II19160));
assign g28651 = ((~g27981));
assign II30044 = ((~g22731));
assign g30981 = ((~II41117));
assign II26567 = (g18679&g14910&g13687);
assign II25300 = (g18708&g18735&g18789);
assign II14037 = ((~g2351));
assign g20325 = ((~g17336));
assign g10313 = (g7015&g1813);
assign g29083 = ((~g28331)&(~g28333));
assign g21194 = (g20250&g12382);
assign g26791 = (g24952&g26525&g13649);
assign II24102 = ((~g6363))|((~g14011));
assign g16449 = (g5985&g12149);
assign g26787 = (g26129&g16636);
assign g9101 = (g3806&g2564);
assign g27889 = ((~II36347));
assign g24447 = ((~g23644))|((~g3306));
assign gbuf37 = (g342);
assign g8270 = ((~II15478));
assign g10509 = (g3494&g1288);
assign g21418 = (g6290&g19705);
assign g15349 = (g4526&g12759);
assign g22497 = ((~II29043));
assign g29991 = (g29901&g8403);
assign g26358 = ((~II34321));
assign g25675 = ((~II33501));
assign g10266 = ((~II17228));
assign g9439 = (g6314&g8126);
assign II33695 = ((~g24538));
assign II35017 = ((~g26616));
assign g22713 = ((~II29395));
assign g23619 = ((~II30735));
assign g6061 = ((~II14562));
assign g19388 = ((~g17139));
assign g10249 = (g3678&g4549);
assign g21960 = ((~II28506));
assign g26607 = ((~g25299)&(~g24578));
assign g22792 = ((~II29562));
assign II25534 = ((~g18179))|((~II25532));
assign g22723 = ((~II29415));
assign g9923 = (g6783&g4159);
assign g30398 = (g30241&g9038);
assign g24803 = (g9795&g24151);
assign II32716 = ((~g23358));
assign g5885 = ((~g2380));
assign II38707 = ((~g29407));
assign II20655 = ((~g12059));
assign g20254 = (g13764&g13797&II26676);
assign g17227 = ((~II23309));
assign II24416 = ((~g14053))|((~II24415));
assign g11636 = ((~II18820));
assign II16009 = ((~g3878));
assign II41019 = ((~g30771))|((~II41017));
assign II39812 = ((~g30312));
assign g6037 = ((~g2273));
assign II28455 = ((~g20943));
assign g15142 = (g4281&g13172);
assign g29551 = ((~II38931));
assign g29160 = ((~II38223));
assign g20395 = ((~II26816));
assign g12017 = ((~g10100));
assign g28378 = (g52&g27776);
assign II33589 = ((~g25069));
assign g10257 = (g7085&g4564);
assign g3948 = ((~g835));
assign g24477 = ((~g24014))|((~g3806));
assign g8853 = ((~II16101));
assign g20444 = ((~g17755));
assign g25346 = (g24644&g18084);
assign g28491 = ((~g27780));
assign g30954 = ((~g30916)&(~g30944));
assign g30259 = ((~g16301)&(~g30093));
assign II25516 = (g17173)|(g17160)|(g17142);
assign g29238 = (g9569&g28814);
assign II23161 = ((~g9453))|((~g13857));
assign II25291 = (g18679&g18699&g18758);
assign g3245 = ((~II13131));
assign g29801 = ((~II39255));
assign II18022 = ((~g6783));
assign II16347 = ((~g5427));
assign g25091 = ((~g23434)&(~g22215));
assign g29341 = (g29062&g29046);
assign g23829 = (g18190&g23038);
assign II37846 = ((~g28501));
assign g13560 = ((~g12711))|((~g3722));
assign g8411 = ((~II15613));
assign g13390 = (g5825&g11459);
assign g28551 = ((~g26038)&(~g27733));
assign II40263 = ((~g30353));
assign II32587 = ((~g17815))|((~II32586));
assign g17197 = ((~g8000)&(~g14259));
assign II25701 = ((~g1435))|((~II25700));
assign g21536 = (g20522)|(g19484)|(g19001);
assign g13269 = ((~II20324));
assign g24845 = ((~g16350)&(~g24246));
assign II36978 = ((~g28053));
assign g28234 = ((~II36951));
assign g25229 = ((~g24777)&(~g23591));
assign g28679 = ((~II37584));
assign g9196 = ((~II16476));
assign g25166 = ((~II32976));
assign gbuf170 = (g2211);
assign g10024 = (g3398&g6912);
assign II14937 = ((~g2003));
assign g9518 = (g3254&g8191);
assign g8805 = ((~II16009));
assign II18347 = ((~g5778));
assign g27539 = ((~II35923));
assign g19452 = ((~g16702));
assign g9145 = (g3774&g7823);
assign II23709 = ((~g13546));
assign g13215 = ((~II20264));
assign g24141 = ((~g22497));
assign g14052 = ((~g11916));
assign II35464 = ((~g26831));
assign g21681 = (g16583&g19534&g14423);
assign g26473 = (g5263&g25838);
assign g21322 = (g9595&g20321);
assign g12451 = ((~g499)&(~g8983));
assign g14273 = ((~g12043));
assign g16558 = (g14863&g14922&g16266&g16360);
assign g13341 = ((~II20414));
assign g16001 = ((~g12601));
assign g22040 = ((~g21307)&(~g19567));
assign g29423 = ((~II38650));
assign II21190 = ((~g13165));
assign II18178 = ((~g6838));
assign II31661 = ((~g23828));
assign g12253 = ((~II19426));
assign g30362 = ((~II39899));
assign g6631 = ((~g2616));
assign g5861 = ((~g930));
assign II18842 = ((~g9084));
assign g21054 = ((~g19903)&(~g18128));
assign g29732 = ((~g6104)&(~g29583)&(~g25387));
assign II37023 = ((~g27799));
assign II35034 = ((~g26087))|((~g26154));
assign II31436 = ((~g22651));
assign II35974 = ((~g27094))|((~g14985));
assign g21398 = (g9277&g20394);
assign g5966 = ((~g1506));
assign II24695 = ((~g6146))|((~II24694));
assign g24174 = ((~g16894)&(~g22206));
assign g24761 = (g9507&g24113);
assign II31024 = ((~g22154));
assign II35482 = ((~g27176));
assign g24797 = ((~II32346))|((~II32347));
assign II29585 = ((~g21045));
assign II17303 = ((~g7391));
assign II33726 = ((~g24557));
assign g12285 = ((~II19455));
assign g12139 = ((~II19318));
assign g12857 = ((~g9326)&(~g9264));
assign g14022 = (g7679&g12921);
assign g8567 = (g3722&g2348);
assign g4392 = ((~g1538));
assign g13209 = ((~g9673));
assign g15461 = ((~II21720));
assign II31144 = ((~g22935));
assign II35859 = ((~g26810));
assign g9885 = ((~g6905));
assign II35422 = ((~g26830));
assign g7912 = ((~g2552));
assign II16283 = ((~g6046));
assign g29969 = (g29721&g22237);
assign g19606 = (g3954&g17360);
assign g10151 = (g3566&g4392);
assign g16501 = ((~g14158));
assign g9066 = (g5512&g7635);
assign g23548 = ((~II30598));
assign g25329 = ((~g24844));
assign II21127 = ((~g12544));
assign II19718 = ((~g8726));
assign g8751 = (g6486&g7906);
assign g5647 = ((~g301));
assign II30158 = ((~g22763));
assign g9498 = ((~II16661));
assign g21112 = (g20250&g12259);
assign II22521 = ((~g13632));
assign g11805 = (g6173&g8643);
assign g20372 = ((~g17476));
assign g29252 = (g28859&g8863);
assign g25787 = ((~II33624));
assign g25154 = ((~II32940));
assign II35976 = ((~g14985))|((~II35974));
assign g13488 = (g6025&g12218);
assign g13115 = ((~g9676))|((~g7162));
assign g4176 = ((~g2079));
assign g27242 = (g26793&g8357);
assign g16184 = (g5663&g11853);
assign g29951 = (g29777&g28945);
assign g24130 = ((~g22480));
assign g21368 = (g9174&g20367);
assign g19145 = ((~II25334));
assign g11173 = ((~II18091));
assign g27195 = ((~II35422));
assign g17174 = ((~g14669))|((~g14691));
assign g13538 = ((~g12565))|((~g3254));
assign II40790 = ((~g30814));
assign II18722 = ((~g8909));
assign g17076 = ((~g14725)&(~g14703)&(~g15923));
assign g24329 = ((~II31661));
assign g5472 = ((~II14006));
assign II37284 = ((~g28147));
assign II22800 = ((~g13581));
assign g15730 = (g5305&g13298);
assign g17430 = ((~II23518));
assign g8007 = ((~II15299));
assign g10381 = (g3522&g4788);
assign g9004 = (g3806&g2571);
assign g26694 = ((~II34689));
assign g15049 = ((~II21404));
assign II22885 = ((~g13370))|((~II22884));
assign g16498 = ((~g14158)&(~g14347));
assign II22803 = ((~g14753));
assign g4581 = ((~g2777));
assign g30408 = ((~II39976));
assign g28650 = ((~g27977));
assign g3566 = ((~II13200));
assign II35993 = ((~g27106))|((~II35992));
assign g6676 = ((~g559));
assign g24221 = (g22979&g11042);
assign g6418 = ((~g1196));
assign g16098 = ((~g12840));
assign g26546 = ((~g25484));
assign II31502 = ((~g23612));
assign g10891 = ((~II17762));
assign g27382 = ((~II35715))|((~II35716));
assign II27281 = ((~g19369));
assign g26678 = ((~II34641));
assign II17780 = ((~g7348));
assign g11718 = ((~g9676))|((~g3522));
assign II36592 = ((~g27529))|((~II36591));
assign g22865 = ((~g16164)&(~g20928));
assign g22257 = ((~g20676));
assign II33327 = ((~g25017));
assign g13481 = (g5864&g11603);
assign II32462 = ((~g24057))|((~II32460));
assign g25219 = ((~g24761)&(~g23572));
assign g16764 = ((~g14976));
assign g26561 = ((~g25524));
assign g20305 = ((~g17291));
assign g22337 = (g2160&g21627);
assign II40847 = ((~g30830));
assign g10004 = ((~II16972));
assign g30274 = ((~g16403)&(~g30108));
assign II19971 = (g9649&g9569&g9453&g9374);
assign II22506 = ((~g13624));
assign g7652 = ((~g1001));
assign g25264 = ((~g24876)&(~g23849));
assign g11823 = ((~g9635)&(~g9763)&(~g9891));
assign g4787 = ((~g1282));
assign g4602 = ((~g525));
assign g10067 = ((~II17027));
assign g10773 = ((~g6431));
assign g19303 = (g16867&g16543&g14071);
assign g28493 = (g18526&g28187);
assign g12608 = ((~II19756));
assign g17262 = ((~II23348));
assign II21803 = ((~g11709));
assign II37303 = ((~g27802))|((~g27900));
assign g10532 = (g7391&g5115);
assign g28188 = (g27349&g11008);
assign g16302 = ((~g13046));
assign II39273 = ((~g29701));
assign g21759 = ((~g20164))|((~g6232));
assign g5361 = ((~g2694));
assign g12117 = ((~g11468));
assign II27379 = ((~g19358));
assign II36301 = ((~g27382))|((~II36300));
assign g16119 = (g3460&g11809);
assign g20943 = ((~II27491));
assign gbuf106 = (g1258);
assign g22659 = ((~II29283));
assign g15764 = ((~g12421));
assign g29558 = (g28790&g29389);
assign g11420 = (g6314&g216);
assign g9770 = ((~II16814));
assign II37991 = ((~g28556));
assign g19448 = ((~g16694));
assign g20377 = ((~II26796));
assign g19037 = ((~II25174));
assign II38196 = ((~g29094));
assign g6209 = ((~g1319));
assign g22253 = ((~II28825));
assign g19234 = (g18578)|(g18611);
assign g25847 = ((~II33689));
assign g13325 = ((~II20394));
assign g13868 = ((~g11633));
assign g29509 = ((~II38857));
assign g23740 = (g17993&g23012);
assign II38071 = ((~g28355));
assign g15139 = ((~II21452));
assign II37029 = ((~g28016));
assign g21382 = ((~II27927));
assign II37566 = ((~g28370));
assign II40039 = ((~g30255));
assign g25928 = ((~g24965))|((~g5438));
assign g20484 = ((~II26931));
assign g18485 = ((~g15756));
assign II34993 = ((~g26575));
assign II23608 = ((~g15889));
assign g10677 = ((~g3398))|((~g6912));
assign g14966 = ((~g11902));
assign g13500 = (g5911&g11633);
assign g28308 = ((~II37173));
assign II17998 = ((~g5668));
assign g7919 = ((~g2963));
assign g5926 = ((~g195));
assign g30883 = ((~II40901));
assign g22197 = ((~II28742))|((~II28743));
assign g18848 = ((~g15308));
assign g16864 = (g15790&g8681);
assign g9110 = (g5556&g7727);
assign g18944 = ((~II24982));
assign g22056 = ((~g21321)&(~g19588));
assign g25798 = ((~g24739)&(~g24526));
assign II36744 = ((~g27333));
assign g17448 = (g4118&g15109);
assign g4234 = ((~g818));
assign II32964 = ((~g24886));
assign g14292 = ((~g12949));
assign g16055 = ((~g12786));
assign g7471 = ((~g3036));
assign g21553 = (g9857&g20476);
assign II33711 = ((~g25073));
assign g18110 = ((~g14107));
assign g26372 = (g4922&g25661);
assign g23918 = ((~g22036));
assign g23147 = ((~g21825));
assign g24273 = ((~II31493));
assign II21449 = ((~g13047));
assign II29339 = ((~g20955));
assign g16368 = (g5915&g12001);
assign g10057 = (g6980&g4260);
assign g17788 = ((~II23863));
assign g5868 = ((~g1609));
assign g22523 = ((~II29073));
assign g27329 = ((~g27081)&(~g26438));
assign II27917 = ((~g19153));
assign g20458 = ((~II26895));
assign II41012 = ((~g30779))|((~II41010));
assign g21902 = ((~g19978));
assign g11091 = ((~II18001));
assign g11797 = ((~g10983));
assign g27704 = ((~II36123));
assign g30892 = ((~II40928));
assign II24531 = ((~g6707))|((~II24530));
assign g23612 = ((~II30722));
assign g20286 = ((~g17249));
assign g18553 = ((~II24625))|((~II24626));
assign II15998 = ((~g3650));
assign II15613 = ((~g7085));
assign g28095 = ((~II36718));
assign g29448 = ((~II38725));
assign II26051 = ((~g16824));
assign g9592 = ((~II16703));
assign g26314 = ((~II34274));
assign II20816 = ((~g12487));
assign g5809 = ((~g780));
assign g22769 = ((~II29525));
assign II34674 = ((~g26211));
assign g12160 = ((~g8357));
assign II18515 = ((~g8843));
assign g11959 = ((~g11249));
assign g30498 = ((~II40086));
assign g7559 = ((~g2565));
assign g25417 = ((~g24830));
assign g18783 = ((~g15034));
assign g8465 = (g6232&g258);
assign g21325 = (g9737&g20324);
assign II30864 = ((~g22493));
assign g6146 = ((~g1358));
assign gbuf160 = (g1862);
assign II36496 = ((~g27267));
assign g14577 = ((~g12234));
assign g27341 = ((~g27097)&(~g26470));
assign g10946 = ((~II17843));
assign g29956 = (g29780&g28998);
assign II33804 = ((~g25976));
assign g30507 = ((~II40101));
assign g18824 = ((~g15185));
assign II16432 = ((~g3366));
assign g29949 = (g29781&g28932);
assign g11549 = ((~II18623));
assign II17875 = ((~g7976));
assign g15902 = (g7607&g2920&II22136);
assign g15639 = (g5216&g13262);
assign g28481 = (g18314&g27981);
assign g15582 = ((~II21838));
assign II17746 = ((~g8107));
assign g12195 = ((~g10437)&(~g10497)&(~g10558));
assign g26807 = ((~g15245)&(~g26261));
assign g14954 = ((~II21351));
assign g26104 = ((~II33999));
assign g26293 = (g4606&g25536);
assign g23144 = ((~g21825));
assign g22786 = ((~II29550));
assign g8548 = (g3410&g888);
assign g10673 = (g7303&g2688);
assign g28624 = ((~g27879));
assign g11733 = ((~g9968))|((~g3834));
assign g19055 = ((~II25228));
assign g21860 = ((~g18270))|((~g19201))|((~g19209));
assign g28219 = ((~II36906));
assign g24097 = ((~g22382));
assign g20417 = ((~g16907)&(~g13833));
assign g4153 = ((~g1413));
assign g13020 = ((~g9534))|((~g6912));
assign g18927 = ((~g15599));
assign g9356 = ((~g5665));
assign g26044 = ((~g25552)&(~g24882));
assign II14609 = ((~g1152));
assign g27994 = ((~II36479));
assign g5636 = ((~g2175));
assign g30347 = ((~II39866));
assign II13107 = ((~g5));
assign g18996 = ((~II25074));
assign II13940 = ((~g1739));
assign g9416 = ((~II16605));
assign g11653 = ((~g9083)&(~g9100)&(~g9109));
assign II34809 = ((~g26249));
assign g11740 = ((~g10877));
assign g26235 = (g25895&g9368);
assign g25324 = ((~II33154));
assign II19634 = ((~g10835));
assign g26782 = ((~II34901));
assign II40910 = ((~g30747));
assign g25238 = ((~g24794)&(~g23611));
assign g15970 = ((~g12711))|((~g6838));
assign g10120 = (g5473&g4372);
assign II17795 = ((~g7976));
assign II20009 = ((~g8313));
assign g30444 = (g30139&g11132);
assign II15859 = ((~g5638));
assign g8103 = ((~g185));
assign g4908 = ((~g734));
assign g30321 = ((~II39806));
assign II15212 = ((~g2947))|((~II15211));
assign gbuf195 = (g2472);
assign g19099 = (g14811&g18699&g18728&g16351);
assign g23526 = ((~g10735))|((~g14584))|((~g22364));
assign g27574 = ((~g26935)&(~g24720));
assign II15876 = ((~g3650));
assign II24015 = ((~g13907))|((~g9427));
assign g29716 = ((~g29498));
assign g13135 = ((~g8626)&(~g8635)&(~g8650));
assign II16104 = ((~g6448));
assign g27300 = ((~g27034)&(~g26372));
assign II31286 = ((~g22267));
assign II40501 = ((~g30682));
assign II39375 = ((~g29768))|((~g15942));
assign g30855 = ((~II40817));
assign g29960 = (g29786&g29050);
assign g9016 = ((~II16338));
assign g27666 = (g26849&g11243);
assign g11228 = ((~II18154));
assign g30605 = ((~g6119)&(~g30412)&(~g25333));
assign g4529 = ((~g1513));
assign g26825 = ((~g15507)&(~g26390));
assign g10693 = (g7462&g7522&g2924&g7545);
assign g24734 = ((~II32248));
assign g19856 = (g4851&g17856);
assign g8696 = ((~II15896));
assign g10539 = (g3834&g5132);
assign g17714 = (g4578&g15376);
assign II30636 = ((~g22037));
assign II14760 = ((~g405));
assign g29211 = (g15210&g28768);
assign g21714 = ((~g20164))|((~g6232));
assign g13845 = (g7559&g12644);
assign g9780 = (g6519&g4041);
assign g17204 = ((~g8075)&(~g14381));
assign g30084 = ((~II39585));
assign g22212 = ((~g21914));
assign g10060 = (g6783&g4269);
assign II27275 = ((~g19369));
assign g28749 = ((~g15064)&(~g28444));
assign g19327 = ((~g14747))|((~g8594))|((~g17130));
assign II21974 = ((~g11726));
assign II32379 = ((~g18247))|((~II32378));
assign g26015 = ((~II33897));
assign g6905 = ((~g3104));
assign II23067 = ((~g14123))|((~II23065));
assign g27153 = ((~g26429));
assign II31547 = ((~g23454));
assign g18645 = (g14776&g14895&g16142&g13750);
assign II21612 = ((~g13062));
assign g13704 = (g7581&g12542);
assign g5798 = (g2400&g2439);
assign g23635 = ((~II30769));
assign II26437 = ((~g16655));
assign g28658 = ((~g27773)&(~g27364));
assign g20608 = ((~II27149));
assign II37232 = ((~g28200));
assign g29180 = (g28982&g20714);
assign II30017 = ((~g22824));
assign g3998 = ((~g23));
assign g29328 = ((~II38505));
assign II16967 = ((~g4452))|((~II16965));
assign g11576 = ((~II18704));
assign g20772 = ((~II27361));
assign II14839 = ((~g2214));
assign g16129 = ((~g12863));
assign g24787 = ((~II32324))|((~II32325));
assign g3975 = ((~g1552));
assign II20706 = ((~g11490));
assign g15574 = ((~II21830));
assign II33286 = ((~g24426));
assign g16849 = ((~II22823));
assign g10683 = ((~g8245));
assign II25938 = ((~g2156))|((~g18142));
assign g27320 = ((~g27062)&(~g26415));
assign g22180 = ((~g21482)&(~g19814));
assign g11495 = ((~II18461));
assign g29635 = ((~II39023));
assign II25717 = ((~g17209));
assign II25791 = ((~g2133))|((~II25790));
assign g4278 = ((~g1561));
assign g5665 = ((~g105));
assign g8907 = (g7078&g5598);
assign II18127 = ((~g6232));
assign g21661 = ((~g19091));
assign g16966 = (g7529&g15174);
assign g24766 = ((~II32285))|((~II32286));
assign g9170 = ((~II16462));
assign g17156 = (g8164&g15738);
assign g30411 = (g30143&g11039);
assign g16719 = ((~II22737));
assign g23723 = (g17954&g23007);
assign II15442 = ((~g3235));
assign g20390 = ((~g17534));
assign II32519 = ((~g18014))|((~II32518));
assign g29106 = ((~II38107));
assign II25032 = ((~g13507))|((~II25030));
assign II16444 = ((~g3678));
assign g30636 = ((~g16140)&(~g30409));
assign g23463 = ((~II30501));
assign g18965 = ((~g15744));
assign g8262 = ((~II15454));
assign g10086 = ((~II17048));
assign g22187 = (g21564&g20986);
assign g21943 = ((~II28455));
assign II36217 = ((~g27580));
assign II14602 = ((~g2530));
assign g17201 = ((~II23278))|((~II23279));
assign g17853 = (g4833&g15496);
assign g6016 = ((~g210));
assign g15789 = ((~g12657))|((~g6783));
assign g29540 = (g26041&g29378);
assign II38360 = ((~g29111));
assign g22317 = ((~g21152))|((~g21241))|((~g21136));
assign II23180 = ((~g9488))|((~II23179));
assign g4049 = ((~g1385));
assign II23103 = ((~g9342))|((~g14052));
assign g29172 = ((~g28846)&(~g28401));
assign II22937 = ((~g9150))|((~II22936));
assign g4171 = ((~g1560));
assign g18140 = (g5196&g15691);
assign II31946 = ((~g23916));
assign g26722 = ((~II34773));
assign II23274 = ((~g13741));
assign g17814 = (g4760&g15467);
assign g12135 = ((~g8324));
assign g8126 = ((~g149));
assign g5707 = ((~g109));
assign g28403 = ((~g27811)&(~g22344));
assign g26387 = (g4997&g25688);
assign g20492 = (g17258&g11894);
assign g19551 = (g16974&g16797&g15003);
assign II18262 = ((~g7195));
assign II16489 = ((~g6000));
assign g13992 = ((~g12836));
assign g18331 = ((~g14626));
assign g21726 = ((~g19105));
assign g9604 = (g6783&g8227);
assign II32423 = ((~g18155))|((~II32422));
assign g29088 = ((~g9507))|((~g28512));
assign g12012 = (g8015&g8745);
assign g19774 = (g1332&g18874);
assign g19320 = (g16867&g16515&g14158);
assign II15971 = ((~g7195));
assign g13181 = ((~g9404));
assign g28048 = ((~II36601));
assign g9648 = (g6678&g3945);
assign II34977 = ((~g26559));
assign g5296 = ((~g1306));
assign g27680 = (g26983&g11392);
assign g23886 = (g18341&g23064);
assign g21565 = ((~g19291));
assign g3925 = ((~g155));
assign g26474 = ((~II34438));
assign II30119 = ((~g22791));
assign g30024 = ((~g29550)&(~g29957));
assign II15204 = ((~g2969))|((~g2972));
assign g9241 = (g6232&g7950);
assign II41047 = ((~g30937));
assign II33643 = ((~g25061));
assign g30489 = (g30175&g11395);
assign g23123 = ((~g17128)&(~g21194));
assign g27108 = (g23395&g26657);
assign g22868 = ((~g21222));
assign II33708 = ((~g24475));
assign II20568 = ((~g13269));
assign g9810 = (g6783&g4067);
assign g10100 = ((~II17070));
assign g19588 = (g8215&g17321);
assign g27415 = ((~g23104)&(~g27181)&(~g25128));
assign g19567 = (g8138&g17282);
assign g30113 = (g29885&g11444);
assign g5702 = ((~g56));
assign II20631 = ((~g11611));
assign II38480 = ((~g28761));
assign g23879 = ((~II31141));
assign g20786 = ((~II27375));
assign g3919 = ((~g3080));
assign g24308 = ((~II31598));
assign g11950 = ((~g11237));
assign g20197 = (g13677&g13706&II26639);
assign g29931 = ((~II39392))|((~II39393));
assign g25615 = ((~II33440));
assign II19791 = ((~g10486));
assign II23917 = ((~g13562));
assign g27305 = ((~g27045)&(~g26383));
assign II22509 = ((~g13610));
assign g27100 = (g23395&g26653);
assign g30977 = ((~II41105));
assign g13438 = ((~II20613));
assign g12495 = ((~g10767));
assign g23942 = (g22980&g10176);
assign II25389 = ((~g18780));
assign g23403 = ((~g23052));
assign g7533 = ((~g1871));
assign II23036 = ((~g13864))|((~II23034));
assign g16005 = ((~g12608));
assign g8515 = (g3254&g192);
assign g17661 = ((~II23745));
assign II35926 = ((~g26821));
assign g27367 = ((~II35689));
assign II29389 = ((~g20974));
assign II16002 = ((~g7391));
assign g11758 = ((~g8514));
assign g8481 = (g3722&g2294);
assign g4112 = ((~g428));
assign g24562 = ((~II32102));
assign g20575 = ((~II27050));
assign g26033 = (g25395&g19452);
assign II36390 = ((~g27243));
assign g6119 = ((~g2574));
assign g23288 = ((~II30317));
assign g11937 = ((~II19119));
assign g15268 = ((~II21551));
assign g25045 = ((~g23955))|((~g6945));
assign g24393 = ((~II31853));
assign II25653 = ((~g1430))|((~g17937));
assign g25892 = ((~g4985)&(~g25099)&(~g18616)&(~g16223));
assign g23006 = ((~g21483));
assign g28775 = ((~II37736));
assign g5961 = ((~g951));
assign g15236 = ((~g12181));
assign g30813 = ((~II40691));
assign g29672 = ((~g29536)&(~g29312));
assign g5413 = ((~II13953));
assign g24013 = ((~g4985)&(~g22997));
assign g16028 = (g5543&g11745);
assign II23763 = ((~g15941));
assign g21389 = (g9649&g20384);
assign II39011 = ((~g29530));
assign g16278 = ((~g12292));
assign g19792 = ((~II26231));
assign g14201 = ((~g11991));
assign II25156 = ((~g18895));
assign g4680 = ((~g1544));
assign g13198 = ((~g9585));
assign g4450 = ((~II13478));
assign g30056 = ((~g29966)&(~g13345));
assign II15457 = ((~g3240));
assign g24933 = ((~g23518));
assign II34746 = ((~g26187));
assign II23745 = ((~g13549));
assign g14336 = (g8099&g12998);
assign g5942 = ((~II14402));
assign g21814 = (g16558)|(g19080)|(g16513)|(II28341);
assign g30835 = ((~II40757));
assign g8947 = (g7328&g5615);
assign II38599 = ((~g29013));
assign g25852 = ((~g4456)&(~g14831)&(~g25078));
assign g29811 = (g29703&g20644);
assign g21969 = ((~g20895)&(~g10133));
assign II13965 = ((~g2433));
assign II17150 = ((~g7465))|((~II17149));
assign II24555 = ((~g14537))|((~II24553));
assign g10569 = (g6751&g1300);
assign II38755 = ((~g29278));
assign II36921 = ((~g28047));
assign g30701 = ((~g13970)&(~g30389));
assign g12559 = ((~g8719));
assign II40239 = ((~g30378));
assign g22058 = ((~g21323)&(~g19590));
assign g25172 = ((~II32994));
assign g20294 = (g18744&g15080&g16433);
assign g22333 = (g21766&g12370);
assign II16179 = ((~g5512));
assign g11862 = ((~g11091));
assign g21537 = ((~II28072));
assign g25436 = ((~II33260));
assign II33849 = ((~g25824));
assign II19689 = ((~g10016));
assign g26497 = ((~g25818));
assign g24127 = ((~g22470));
assign II31922 = ((~g23543));
assign g24354 = ((~II31736));
assign g14922 = ((~g12214));
assign II15398 = ((~g2845));
assign g13305 = ((~g8317))|((~g2993));
assign II21064 = ((~g13147));
assign g22185 = ((~g21490)&(~g19824));
assign II30467 = ((~g23000));
assign g25191 = ((~g24516)&(~g22777));
assign g15172 = (g4346&g13176);
assign g4111 = ((~g420));
assign II39457 = ((~g29943));
assign g8487 = (g6232&g267);
assign II33703 = ((~g24545));
assign g16026 = ((~g12708));
assign g17410 = ((~II23498));
assign g19053 = ((~II25222));
assign g7555 = ((~g1152));
assign g15112 = ((~II21432));
assign II13211 = ((~g1930));
assign g15265 = ((~II21548));
assign g6034 = ((~g1588));
assign g21770 = ((~g14490))|((~g15355))|((~g19927))|((~g19906));
assign g7570 = ((~g3032));
assign g23406 = ((~g17597)&(~g22618));
assign g7658 = ((~g1090));
assign II27059 = ((~g19207));
assign II25914 = ((~g1462))|((~II25913));
assign g28235 = ((~II36954));
assign II34743 = ((~g26118));
assign g20531 = ((~II26972));
assign g25817 = ((~II33655));
assign g24433 = (g24134&g13626);
assign g13978 = ((~g11873));
assign g24248 = ((~II31436));
assign g9621 = (g7085&g8236);
assign g8278 = ((~g3337));
assign II30287 = ((~g22692));
assign g8946 = (g7303&g2565);
assign g21967 = ((~II28527));
assign g29232 = (g9356&g28796);
assign g28112 = (g27622&g10266);
assign g27492 = ((~g24958)&(~g24633)&(~g26771));
assign g26728 = ((~II34791));
assign II17632 = ((~g6183));
assign g10940 = ((~II17837));
assign II30248 = ((~g22599));
assign II27080 = ((~g19198));
assign g23047 = ((~g16991)&(~g21103));
assign g9338 = ((~II16559));
assign g28092 = ((~II36711));
assign II36984 = ((~g28013));
assign g26788 = ((~II34909));
assign II37605 = ((~g28583));
assign g19876 = (g17842&g18297&II26320);
assign g30476 = (g30175&g11318);
assign g18538 = ((~II24602))|((~II24603));
assign g8084 = ((~g2563));
assign g25048 = ((~g23984))|((~g7053));
assign g14337 = ((~II21165));
assign g27915 = (g13936&g27410);
assign g17812 = (g4754&g15461);
assign g16399 = ((~II22444));
assign g30532 = ((~II40176));
assign g20491 = ((~II26940));
assign g26603 = ((~g25655));
assign g15231 = ((~II21514));
assign g23718 = ((~II30888));
assign g30458 = (g30159&g11219);
assign g26540 = ((~g25467));
assign g8801 = (g3806&g8164);
assign II38680 = ((~g29404));
assign g21090 = ((~g19064));
assign g21124 = (g19471&g18004&g14194);
assign g10310 = (g3566&g4680);
assign g8468 = (g6369&g936);
assign g30772 = ((~II40578));
assign II37266 = ((~g28200));
assign g5778 = ((~g1680));
assign g5968 = ((~g1636));
assign g8904 = ((~II16182));
assign g9606 = (g6574&g8233);
assign g27301 = ((~g27035)&(~g26373));
assign II23772 = ((~g15055));
assign II25186 = ((~g18998));
assign II27534 = ((~g20083));
assign g30791 = ((~II40628))|((~II40629));
assign g23028 = ((~g21541));
assign II23154 = ((~g14061))|((~II23152));
assign g9901 = (g3366&g4115);
assign gbuf10 = (g2830);
assign II14069 = ((~g1564));
assign II23545 = ((~g15867));
assign g18358 = ((~g14360));
assign g5283 = ((~g2795));
assign g28436 = (g17954&g28161);
assign g8941 = ((~II16241));
assign g30939 = ((~II41041));
assign II28346 = (g20277)|(g20268)|(g20247);
assign g28190 = ((~g27555));
assign g29103 = ((~g9795))|((~g28567));
assign II38548 = ((~g28903));
assign g27809 = ((~II36271))|((~II36272));
assign g4897 = ((~g602));
assign II28984 = ((~g21747));
assign g9184 = ((~II16472));
assign g22178 = ((~g21480)&(~g19812));
assign g23280 = ((~II30293));
assign g13113 = ((~g9534))|((~g6912));
assign II16332 = ((~g3462));
assign g22063 = ((~g21328)&(~g19597));
assign g16186 = (g5753&g11856);
assign II38363 = ((~g29016));
assign g22741 = ((~II29459));
assign g25873 = ((~g4632)&(~g14904)&(~g25082));
assign g13326 = (g2373&g11256);
assign g11259 = ((~II18187));
assign II21726 = ((~g13112));
assign g23468 = ((~II30508));
assign g24059 = ((~g21990)&(~g20809));
assign g24538 = ((~g15581)&(~g23900));
assign II30954 = ((~g14309))|((~II30952));
assign g29386 = ((~g29010));
assign g8717 = (g3338&g7953);
assign g10877 = ((~II17740));
assign II18743 = ((~g9025));
assign II35702 = ((~g26867))|((~II35701));
assign II19924 = ((~g10726));
assign g29542 = ((~II38916));
assign g6890 = ((~g2714));
assign g9809 = (g3566&g4064);
assign II36731 = ((~g27567))|((~g15055));
assign g29921 = ((~g29736)&(~g22367));
assign II23418 = ((~g15824));
assign g25605 = ((~g25096)&(~g6184));
assign g11545 = ((~II18611));
assign g10872 = ((~g5884)&(~g5920)&(~g5949));
assign II37116 = ((~g28068));
assign II25386 = ((~g18763));
assign g27283 = ((~g27017)&(~g26333));
assign g26684 = ((~II34659));
assign g15876 = ((~II22120));
assign g27530 = (g23945&g27153);
assign g16913 = ((~g13589));
assign g26646 = ((~g25811));
assign g3922 = ((~g150));
assign g24340 = ((~II31694));
assign g30445 = (g30147&g11135);
assign II27089 = ((~g20105));
assign II36291 = ((~g15923))|((~II36289));
assign II25889 = ((~g1457))|((~II25888));
assign g27685 = ((~II36066));
assign II17866 = ((~g6713));
assign II33840 = ((~g25779));
assign g26655 = ((~g25328)&(~g17084));
assign g12874 = ((~g8915));
assign II30489 = ((~g22911));
assign g4150 = ((~g1388));
assign g16910 = ((~II22875));
assign g20413 = ((~g17613));
assign g9962 = ((~II16958));
assign g30328 = ((~II39825));
assign g11980 = ((~g10115)&(~g10204)&(~g10291));
assign g10778 = (g2929)|(g8022);
assign g16387 = (g5934&g12038);
assign II30227 = ((~g22832));
assign g26507 = ((~II34479));
assign II36257 = ((~g27527))|((~II36256));
assign g28836 = (g5810&g28491);
assign g17055 = (g7153&g15524);
assign g26721 = ((~II34770));
assign II36593 = ((~g14885))|((~II36591));
assign g11472 = ((~II18438));
assign II30170 = ((~g22626));
assign g27800 = ((~II36253));
assign g19631 = (g4032&g17402);
assign g20571 = ((~II27038));
assign g30273 = ((~g16393)&(~g30107));
assign II40826 = ((~g30810));
assign g13866 = ((~g11772));
assign g19868 = (g16498&g16867&g19001);
assign g16844 = ((~g15754)&(~g12989));
assign II28369 = (g20291)|(g18666)|(g18653);
assign g21119 = ((~g20092)&(~g20115)&(~g20139));
assign g5318 = ((~g2682));
assign g22194 = ((~g21523)&(~g19858));
assign g27107 = (g5266&g26474);
assign II23701 = ((~g15055));
assign g20822 = ((~II27411));
assign g14490 = ((~g12172));
assign g26091 = (g2142&g25860);
assign g16496 = ((~II22590));
assign g16174 = ((~g12952))|((~g2013));
assign II33906 = ((~g25519));
assign g15258 = (g4515&g13188);
assign g12116 = ((~g11465));
assign g11818 = ((~g11011));
assign II40158 = ((~g30376));
assign g18904 = ((~g15513));
assign g29145 = ((~II38178));
assign II20448 = ((~g9050));
assign g29710 = ((~g6104)&(~g29583)&(~g25412));
assign g9665 = (g6369&g3963);
assign II34238 = ((~g25251));
assign g28380 = (g1430&g28014);
assign II32109 = ((~g24206));
assign g15854 = ((~g13353))|((~g12392));
assign g25126 = ((~g24030));
assign g29820 = (g29717&g20743);
assign g9276 = ((~II16524));
assign g12934 = ((~g8974));
assign g22756 = ((~II29490));
assign g24376 = ((~II31802));
assign gbuf89 = (g1044);
assign g28318 = ((~II37203));
assign g5135 = ((~g2807));
assign g15040 = ((~II21395));
assign g20880 = ((~g19602)&(~g17397));
assign II40297 = ((~g30482));
assign g4899 = ((~g716));
assign g29963 = (g29758&g13737);
assign g21327 = ((~II27868));
assign II19621 = ((~g10851));
assign g18786 = ((~g15043));
assign g22161 = ((~g21428)&(~g19764));
assign II32042 = ((~g23399));
assign II34102 = ((~g25220));
assign g21928 = ((~II28443));
assign g12330 = (g8246&g8879);
assign II18533 = ((~g10967));
assign II36290 = ((~g27565))|((~II36289));
assign g11575 = ((~II18701));
assign g13562 = ((~g12711))|((~g3722));
assign g22971 = ((~g21779));
assign II31916 = ((~g23485));
assign II21939 = ((~g13142));
assign II26369 = ((~g17059));
assign g21072 = ((~g19926)&(~g18223));
assign g27340 = ((~g27096)&(~g26469));
assign II24104 = ((~g14011))|((~II24102));
assign g25321 = (g25075&g9669);
assign g17839 = ((~II23904));
assign g16850 = (g6226&g14764);
assign g4717 = ((~g2429));
assign g24132 = ((~g22487));
assign II15288 = ((~g3109));
assign g4127 = ((~g841));
assign g28625 = ((~g28100));
assign g19275 = (g16867)|(g16515)|(g19001);
assign g18257 = ((~II24252))|((~II24253));
assign g17428 = (g3994&g16007);
assign g5947 = ((~g2318));
assign g5946 = ((~g2312));
assign g29683 = ((~g29559)&(~g29337));
assign II30080 = ((~g22649));
assign g10125 = ((~II17097));
assign II39881 = ((~g30283));
assign II20744 = ((~g11621))|((~II20743));
assign g14102 = ((~g11946));
assign g18925 = ((~g15588));
assign g11331 = ((~II18288))|((~II18289));
assign g6086 = ((~II14605));
assign g27939 = ((~II36404));
assign g14642 = ((~II21246));
assign g11117 = ((~II18031));
assign g30845 = ((~II40787));
assign g29060 = ((~g9277))|((~g28595));
assign g3990 = ((~g2245));
assign g19858 = (g4857&g17862);
assign II16593 = ((~g6059));
assign g11829 = ((~g11035));
assign g22903 = ((~II29700));
assign g12748 = ((~g8823));
assign g18164 = (g5230&g15711);
assign II16627 = ((~g6448));
assign II25728 = ((~g17118));
assign g28311 = ((~II37182));
assign g4925 = ((~g1268));
assign II32378 = ((~g18247))|((~g24027));
assign II16766 = ((~g6751));
assign II36078 = ((~g27508));
assign g21944 = ((~II28458));
assign II18581 = ((~g8964));
assign g24594 = ((~II32170));
assign II32937 = ((~g24544));
assign g17753 = (g4659&g15415);
assign g29195 = ((~g28880)&(~g28438));
assign g22966 = ((~g21730));
assign g14774 = ((~II21310));
assign g29349 = ((~II38536));
assign II32910 = ((~g24576));
assign g26656 = ((~g25856));
assign g27205 = ((~II35452));
assign g18993 = ((~II25067));
assign g16455 = (g5991&g12159);
assign g29652 = ((~II39074));
assign g8044 = ((~g3194));
assign g27932 = ((~II36397));
assign g18102 = ((~g14668))|((~g9782));
assign II15803 = ((~g8107));
assign g29938 = ((~II39414));
assign g11284 = ((~II18232));
assign II31085 = ((~g22171));
assign II14449 = ((~g3224));
assign II27646 = ((~g20507));
assign g5512 = ((~II14020));
assign II30601 = ((~g22028));
assign g22122 = ((~g21378)&(~g19692));
assign g21018 = ((~g19849)&(~g15556));
assign g22031 = ((~g21299)&(~g19558));
assign g28899 = ((~II37868));
assign g20537 = ((~g18626))|((~g3036));
assign II13165 = ((~g401));
assign g23039 = ((~g16989)&(~g21098));
assign g25999 = ((~II33849));
assign II38758 = ((~g29279));
assign II40597 = ((~g30706));
assign g9868 = (g3722&g4073);
assign g21108 = ((~II27667));
assign g11954 = ((~g11243));
assign g27049 = (g23353&g26615);
assign II38842 = ((~g29333))|((~II38841));
assign II25595 = ((~g61))|((~g18074));
assign g11032 = ((~II17945));
assign II15211 = ((~g2947))|((~g2953));
assign g23061 = ((~g21793)&(~g21163));
assign g25116 = ((~g23882));
assign II15556 = ((~g6783));
assign g13462 = ((~II20685));
assign g24622 = ((~g23616)&(~g22546));
assign g23909 = (g18453&g23082);
assign g19625 = (g4006&g17390);
assign g15412 = ((~II21674));
assign II34313 = ((~g25265));
assign g26298 = (g4641&g25540);
assign II23725 = ((~g13547));
assign II38163 = ((~g29075));
assign g20917 = ((~g19676)&(~g17544));
assign g26909 = ((~II35106));
assign g22356 = ((~g20813));
assign g20183 = (g14811&g18699&g16201&g16254);
assign g30316 = ((~II39791));
assign II20429 = ((~g11262))|((~g11188));
assign g26626 = ((~g25732));
assign g16380 = (g5925&g12020);
assign g11633 = ((~II18817));
assign g12184 = ((~g10414)&(~g10476)&(~g10536));
assign II32518 = ((~g18014))|((~g24071));
assign g19797 = (g2720&g18882);
assign II25862 = ((~g17177));
assign g23528 = ((~g22936)&(~g5659));
assign II24577 = ((~g14614))|((~II24575));
assign g30558 = ((~II40254));
assign g12208 = ((~g10448)&(~g10512)&(~g10570));
assign g26102 = ((~II33995));
assign g19544 = (g16913&g16728&g14849);
assign g9225 = ((~II16493));
assign II39065 = ((~g29514));
assign g11938 = ((~g10037)&(~g10113)&(~g10201));
assign g11953 = ((~g10066)&(~g10157)&(~g10227));
assign II30973 = ((~g22141));
assign II23833 = ((~g15921));
assign g17985 = ((~g14641))|((~g9636));
assign g26401 = ((~II34363));
assign g5906 = ((~g1496));
assign II31523 = ((~g23642));
assign II24264 = ((~g14342))|((~II24263));
assign g21530 = ((~II28065));
assign g10222 = (g6574&g4532);
assign g27093 = (g22108&g26648);
assign g19590 = (g8227&g17327);
assign g22252 = ((~g20669));
assign g10081 = (g6838&g4310);
assign II24017 = ((~g9427))|((~II24015));
assign II13316 = ((~g2836));
assign II23279 = ((~g14320))|((~II23277));
assign II32883 = ((~g24592));
assign II23510 = ((~g15827));
assign g15446 = ((~II21708));
assign g19934 = ((~II26388));
assign II27250 = ((~g19390));
assign g8227 = ((~g1528));
assign g12535 = ((~g8296))|((~g5512));
assign g23659 = (g22784&g17500);
assign II33990 = ((~g25870));
assign II23655 = ((~g14831));
assign g17767 = ((~II23842));
assign g4249 = ((~g1101));
assign II34453 = ((~g25279));
assign g9374 = ((~g5761));
assign g24274 = ((~II31496));
assign II18151 = ((~g5720));
assign g20212 = ((~g16848));
assign g13484 = (g6021&g12210);
assign II13430 = ((~g101));
assign g11613 = ((~II18791));
assign g23577 = (g3957&g22455);
assign gbuf82 = (g971);
assign g20743 = ((~II27332));
assign II23018 = ((~g9216))|((~g14032));
assign II24726 = ((~g6222))|((~II24725));
assign g15352 = ((~g12253));
assign g24096 = ((~g22405));
assign g10527 = (g3774&g5104);
assign g8206 = ((~g175));
assign g6225 = ((~II14704));
assign g21810 = (g20185)|(g20149)|(II28335);
assign g13505 = (g6039&g12267);
assign g20627 = ((~II27206));
assign g5820 = ((~g1486));
assign g13963 = ((~g12820));
assign g18847 = ((~g15293));
assign g28208 = ((~II36873));
assign II29294 = ((~g20941));
assign g17181 = (g7751&g14329);
assign g10279 = (g3306&g4592);
assign g11163 = ((~II18079));
assign g4468 = ((~g358));
assign g27244 = (g26914&g22258);
assign g5038 = ((~g724));
assign g17967 = (g5015&g15588);
assign II16360 = ((~g7265));
assign g4508 = ((~II13504));
assign g28415 = ((~II37357))|((~II37358));
assign g27193 = ((~II35416));
assign g16855 = (g15722&g8646);
assign g26034 = (g25405&g19479);
assign g18154 = (g5224&g15707);
assign II17278 = ((~g3650));
assign II23487 = ((~g13511));
assign g21178 = (g19524&g14546);
assign II31232 = ((~g22026));
assign g13271 = ((~II20328));
assign g30916 = (g30785&g22251);
assign g19306 = ((~g14719))|((~g8587))|((~g17092));
assign g24298 = ((~II31568));
assign II38202 = ((~g29104));
assign g21602 = (g17937&g18379&g19876&II28133);
assign g26520 = ((~g25874));
assign g30926 = ((~II41011))|((~II41012));
assign g15933 = ((~g11663));
assign II33460 = ((~g24452));
assign II39533 = ((~g29915))|((~II39532));
assign II31865 = ((~g23678));
assign II17557 = ((~g3900));
assign II14034 = ((~g1186));
assign g17353 = (g3945&g14963);
assign II19750 = ((~g8726));
assign g28207 = ((~II36870));
assign g10972 = ((~II17869));
assign g12643 = ((~g8775));
assign g7143 = ((~g2998));
assign II35313 = ((~g26534));
assign g13164 = ((~g8706)&(~g8724)&(~g8760));
assign g19216 = (g18606)|(g18053);
assign g11697 = ((~g9125)&(~g9131)&(~g9133));
assign g21148 = ((~g20138)&(~g20161)&(~g20190));
assign g11491 = ((~II18449));
assign g10152 = (g6783&g4395);
assign g25005 = ((~g23539))|((~g2142));
assign II32150 = ((~g24222));
assign g21518 = ((~II28051));
assign g21741 = ((~g20198))|((~g6519));
assign g22256 = ((~g20673));
assign II14532 = ((~g354));
assign g26837 = ((~II34980));
assign g7593 = ((~g2571));
assign II37768 = ((~g28540));
assign II25249 = ((~g17300));
assign g20119 = (g13714&g13756&II26567);
assign II29073 = ((~g21761));
assign g23913 = ((~g23061)&(~g18636)&(~g4985));
assign g25017 = ((~g23644))|((~g5438));
assign II38811 = ((~g29303))|((~II38810));
assign g20588 = ((~II27089));
assign II31679 = ((~g23453));
assign g10384 = (g3522&g4797);
assign II15863 = ((~g3806));
assign g28682 = ((~II37593));
assign g22440 = ((~II28984));
assign g23772 = (g21825&g22875);
assign g21304 = (g9293&g20296);
assign g13185 = ((~g9443));
assign g16164 = ((~g11953));
assign g19503 = (g16884)|(g16697)|(g16665);
assign g20328 = ((~g17345));
assign II25207 = ((~g16559));
assign g29250 = ((~II38355));
assign II23507 = ((~g13514));
assign II17225 = ((~g7391));
assign g11820 = ((~g11017));
assign II14565 = ((~g461));
assign g8891 = ((~II16159));
assign g23441 = ((~g23129));
assign g11764 = ((~g10921));
assign II23200 = ((~g14176))|((~II23198));
assign g30602 = ((~g6119)&(~g30412)&(~g25417));
assign g4824 = ((~g1765));
assign g11931 = ((~g11205));
assign g19501 = ((~II25939))|((~II25940));
assign g29941 = ((~g16182)&(~g29793));
assign II18764 = ((~g9879));
assign g13210 = ((~g9727));
assign g18556 = ((~II24640))|((~II24641));
assign g10545 = ((~II17486));
assign g28496 = ((~g27787));
assign g23676 = ((~II30826));
assign II34961 = ((~g26545));
assign g30628 = ((~g30412)&(~g2610));
assign II40802 = ((~g30730));
assign g23724 = (g22940&g20438);
assign g19957 = ((~II26413));
assign g24384 = ((~II31826));
assign g29805 = ((~II39267));
assign g30889 = ((~II40919));
assign g7461 = ((~g2175));
assign g29699 = ((~II39151));
assign II25216 = ((~g18999));
assign g17534 = ((~II23622));
assign g20479 = ((~II26926));
assign II24765 = ((~g14573))|((~II24763));
assign g25024 = ((~g23748))|((~g5512));
assign g29342 = (g29107&g29054);
assign II24401 = ((~g9264))|((~II24399));
assign II28450 = ((~g19390));
assign g7390 = ((~II14981));
assign g16325 = ((~g13107));
assign g20051 = (g18063&g3114);
assign g28470 = ((~g27671)&(~g28193));
assign II13125 = ((~g23));
assign g9876 = ((~II16870));
assign g29739 = ((~g29505));
assign II18698 = ((~g11255));
assign g20394 = ((~g17551));
assign g8565 = (g7085&g2273);
assign g19918 = ((~g18646));
assign g26028 = (g25438&g24941);
assign g12136 = ((~II19315));
assign g17658 = ((~II23742));
assign g22867 = ((~II29663));
assign g28453 = (g28137&g9335);
assign g16093 = ((~g12833));
assign g12604 = ((~II19750));
assign g30110 = (g29881&g11417);
assign g27787 = ((~II36230));
assign g14955 = ((~II21354));
assign g29428 = ((~II38665));
assign g23259 = ((~II30230));
assign g12068 = ((~g10271)&(~g10352)&(~g10412));
assign g23113 = ((~g21198)&(~g19385)&(~g19413));
assign II30891 = ((~g22116));
assign g25196 = (g24672&g16640);
assign g10692 = (g3834&g5343);
assign g26785 = ((~g26410))|((~g3618));
assign g5650 = (g325&g364);
assign II37790 = ((~g28595));
assign g20082 = ((~II26512));
assign g17225 = ((~g16008)&(~g16015));
assign II17149 = ((~g7465))|((~g7142));
assign g20102 = (g18053)|(g18606)|(II26538);
assign g19600 = (g633&g18783);
assign g13202 = ((~g9610));
assign g22520 = ((~II29070));
assign g17876 = (g4876&g15516);
assign II20858 = ((~g12539));
assign II25021 = ((~g14546));
assign II23082 = ((~g9310))|((~g13879));
assign II14641 = ((~g2540));
assign g30737 = ((~II40495));
assign g25244 = ((~g24804)&(~g23632));
assign g5405 = ((~II13931));
assign g23856 = ((~II31102));
assign II17048 = ((~g6117));
assign g30706 = ((~g14113)&(~g30394));
assign g5630 = (g325&g349);
assign II31850 = ((~g23634));
assign II25102 = ((~g18944));
assign g26993 = (g21976&g26561);
assign g4404 = ((~g1795));
assign g21707 = (g2892&g19978);
assign II32296 = ((~g18014))|((~II32295));
assign g29554 = ((~II38936));
assign g17268 = (g8024&g15991);
assign g24652 = ((~g24183)&(~g531));
assign g26564 = ((~g25533));
assign g29444 = ((~II38713));
assign g17285 = ((~II23371));
assign II19503 = ((~g10486));
assign g23545 = ((~g22984)&(~g20285));
assign g26707 = ((~II34728));
assign g30251 = ((~g16198)&(~g30085));
assign g19776 = (g1358&g18876);
assign II41096 = ((~g30963));
assign II14094 = ((~g2258));
assign g26237 = ((~g25306));
assign g6064 = ((~II14571));
assign g21153 = (g20054&g16543&g16501);
assign g16437 = ((~II22475));
assign g11857 = ((~g11082));
assign g10052 = ((~II17012));
assign g17815 = ((~II23888));
assign g16403 = (g5948&g12065);
assign g15136 = ((~II21449));
assign g4873 = ((~g2783));
assign g16567 = ((~g15904)&(~g15880)&(~g15859));
assign g21364 = ((~g20486)&(~g13266));
assign II32710 = ((~g14402))|((~II32708));
assign g29239 = (g9595&g28817);
assign g3945 = ((~g726));
assign II18548 = ((~g8792));
assign g17588 = ((~II23676));
assign g11616 = ((~II18794));
assign II30209 = ((~g22765));
assign II30985 = ((~g22992));
assign g29022 = (g14502&g28655);
assign g25070 = ((~g24014))|((~g7391));
assign g13507 = ((~II20744))|((~II20745));
assign II22866 = ((~g13612));
assign g23824 = (g22949&g9641);
assign g22567 = ((~II29129));
assign g20707 = ((~g20198))|((~g3410));
assign g24802 = (g9711&g24150);
assign II27270 = ((~g19335));
assign g14596 = ((~g13022));
assign g17030 = ((~II23009))|((~II23010));
assign g8446 = (g3566&g1600);
assign II26843 = ((~g17228));
assign g25213 = ((~g24752)&(~g23560));
assign g29188 = (g29083&g20796);
assign g9404 = ((~II16601));
assign g21495 = ((~II28031));
assign g18572 = ((~g14558));
assign g15408 = ((~g12282));
assign g29664 = ((~g29552));
assign g13430 = ((~II20589));
assign g4048 = ((~g1142));
assign g27879 = ((~II36341));
assign g21395 = (g15274&g20391);
assign g30750 = (g30593&g20729);
assign g23613 = ((~II30725));
assign g29318 = ((~II38483));
assign g25268 = ((~g24888)&(~g17950));
assign g5882 = (g2412&g2443);
assign II31021 = ((~g22153));
assign g13003 = ((~g9058));
assign g5712 = ((~g305));
assign II29098 = ((~g20879));
assign g11869 = ((~g11102));
assign II29101 = ((~g20880));
assign g21277 = (g19681&g15161);
assign g21766 = ((~g19934));
assign II17689 = ((~g6635));
assign g5138 = ((~g2809));
assign g11114 = ((~II18028));
assign g23779 = ((~II30985));
assign II21178 = ((~g11749));
assign g16560 = ((~g14423));
assign II23406 = ((~g15787));
assign g8501 = (g6232&g195);
assign g5747 = ((~II14191));
assign g14044 = ((~g11914));
assign g22794 = ((~II29566));
assign g19039 = ((~II25180));
assign g18840 = ((~g15254));
assign g21981 = ((~g21254)&(~g21267));
assign II30611 = ((~g22030));
assign g19569 = (g8144&g17288);
assign g25301 = ((~g24952));
assign II33974 = ((~g25389));
assign II23996 = ((~g14337));
assign II40952 = ((~g30727));
assign g29773 = ((~g29474)&(~g29208));
assign g29567 = (g29231&g29396);
assign g23615 = (g4107&g22512);
assign II22548 = ((~g14718));
assign g18593 = ((~g15831));
assign g24404 = ((~II31886));
assign g25169 = ((~II32985));
assign II29472 = ((~g21004));
assign g5864 = ((~g1195));
assign g18131 = ((~II24144));
assign g28330 = (g27864&g20711);
assign g29166 = ((~II38241));
assign g27708 = ((~II36135));
assign g16968 = (g6672&g15176);
assign g16697 = ((~g14837));
assign g8540 = (g3566&g1645);
assign g29451 = ((~II38734));
assign g5395 = ((~II13901));
assign g12909 = ((~g10904));
assign II17901 = ((~g6369));
assign II24327 = ((~g9857))|((~II24325));
assign g5689 = ((~g1444));
assign g17640 = ((~g13873));
assign g25188 = (g24652&g20763);
assign II24669 = ((~g9737))|((~II24667));
assign g28257 = ((~II37020));
assign g17474 = (g4176&g15145);
assign g28664 = (g27997&g12055);
assign g13983 = ((~g12828));
assign II29852 = ((~g21331));
assign g20939 = ((~g19722)&(~g17632));
assign g27198 = ((~II35431));
assign g12992 = ((~g8539)&(~g8552)&(~g8561));
assign g25043 = ((~g23694))|((~g5473));
assign g10977 = ((~II17878));
assign g28328 = ((~g27755)&(~g10340));
assign g29108 = ((~II38111));
assign g24978 = (g23954)|(g23974);
assign g23865 = (g22966&g9816);
assign g14032 = ((~g11906));
assign g29673 = ((~g29583));
assign II28314 = ((~g19152));
assign g11358 = ((~II18314));
assign g20569 = ((~II27032));
assign g19814 = (g4680&g17761);
assign g14668 = ((~g11865));
assign II33995 = ((~g25935));
assign g12449 = ((~II19621));
assign II37053 = ((~g28062));
assign g30272 = ((~g16392)&(~g30106));
assign II14769 = ((~g545));
assign g11586 = ((~II18734));
assign g30789 = ((~g30575)&(~g22387));
assign g23877 = (g18314&g23060);
assign g19176 = ((~II25389));
assign g26389 = (g25264&g17962);
assign g28260 = ((~II37029));
assign II40559 = ((~g30605))|((~II40558));
assign gbuf108 = (g1252);
assign g11716 = ((~g9534))|((~g3366));
assign g18967 = ((~g15750));
assign g28802 = ((~g28492)&(~g28036));
assign g4044 = ((~g866));
assign g5984 = ((~g885));
assign g20131 = (g18486&g3176);
assign II35681 = ((~g26869));
assign g27713 = ((~II36150));
assign g12086 = ((~g11432));
assign g27117 = ((~g26320))|((~g6448));
assign g4574 = ((~g2495));
assign g19926 = (g2066&g18963);
assign g14256 = ((~g12036));
assign II16141 = ((~g5409));
assign g23194 = ((~II30035));
assign g9124 = (g6448&g7769);
assign II21790 = ((~g13099));
assign II35434 = ((~g27150));
assign II18820 = ((~g10890));
assign g28683 = ((~II37596));
assign g18972 = ((~g15766));
assign g21848 = ((~g17807))|((~g19181))|((~g19186));
assign gbuf72 = (g823);
assign g24683 = (g17214&g24153);
assign g23424 = ((~g23100));
assign g23349 = ((~g23029))|((~g22198));
assign g11660 = ((~g8183)&(~g8045)&(~g7928)&(~g11069));
assign g9595 = ((~g5775));
assign g7603 = ((~g3133));
assign g7482 = ((~g1842));
assign II14816 = ((~g1092));
assign II37623 = ((~g28467));
assign II30560 = ((~g23110));
assign II28096 = (g13907&g14238&g13946);
assign g24216 = ((~g16994)&(~g22255));
assign g25376 = ((~g24852));
assign II27343 = ((~g19431));
assign II31604 = ((~g23575));
assign g15460 = (g4898&g13219);
assign g24231 = ((~g17048)&(~g22292));
assign g23889 = (g22962&g9913);
assign g27659 = (g27132&g11114);
assign g13885 = ((~g11799));
assign g18879 = ((~g15432));
assign g19709 = (g1339&g18842);
assign g19954 = ((~g17186))|((~g92));
assign g16665 = ((~g14776));
assign g29213 = ((~g15235)&(~g28949));
assign g18400 = ((~g14420));
assign g5693 = ((~g1506));
assign II23564 = ((~g13526));
assign g11992 = ((~g10150)&(~g10221)&(~g10308));
assign II40964 = ((~g30753));
assign II25625 = ((~g18374))|((~II25623));
assign g30731 = ((~II40481));
assign g27725 = (g27532&g20704);
assign II29064 = ((~g20875));
assign g7972 = ((~g3059));
assign II37823 = ((~g28384))|((~II37822));
assign g19236 = (g16935&g8802);
assign II34195 = ((~g25244));
assign g23686 = (g17882&g22998);
assign g17190 = ((~II23257))|((~II23258));
assign g29135 = ((~II38148));
assign g19586 = (g8209&g17315);
assign gbuf183 = (g2365);
assign II19847 = ((~g10677));
assign II22022 = ((~g13145));
assign g24458 = ((~g23694))|((~g3462));
assign g9095 = (g5473&g7682);
assign II31550 = ((~g23481));
assign II18046 = ((~g3254));
assign g8418 = ((~II15620));
assign g20558 = ((~II26999));
assign g28881 = (g28612&g9199);
assign g18809 = ((~g15130));
assign g13102 = ((~g9676))|((~g6980));
assign II27395 = ((~g19431));
assign II24611 = ((~g15814))|((~g15978));
assign g10440 = (g6713&g4916);
assign g10507 = (g6945&g5050);
assign g4343 = ((~g369));
assign g19784 = (g2033&g18877);
assign II17238 = ((~g3900));
assign g18981 = ((~II25037));
assign g20553 = ((~g18569));
assign g28595 = (g26520)|(g27756);
assign g24167 = ((~g22573));
assign II32393 = ((~g24034))|((~II32391));
assign g5875 = ((~g2124));
assign g18236 = ((~g14230));
assign II30290 = ((~g22663));
assign g10194 = (g6448&g4468);
assign g21349 = (g9248&g20347);
assign g10536 = (g3834&g5123);
assign g3833 = ((~g2574));
assign g12169 = ((~g10394)&(~g10456)&(~g10517));
assign g19047 = ((~II25204));
assign g29269 = ((~g28755));
assign g13945 = ((~g11855));
assign gbuf155 = (g1952);
assign g11557 = ((~II18647));
assign g7227 = ((~g1839));
assign g20006 = (g5358&g18466);
assign gbuf171 = (g2256);
assign g29526 = (g27741&g29367);
assign II22590 = ((~g13863));
assign g11844 = ((~g9748)&(~g9871)&(~g9955));
assign g30356 = ((~g14419)&(~g30227));
assign g30076 = ((~II39573));
assign g24759 = (g21825&g23885);
assign g17620 = (g4418&g15293);
assign g17545 = ((~II23633));
assign II38719 = ((~g29258));
assign g27952 = ((~II36417));
assign g11306 = ((~II18256));
assign g28697 = ((~II37638));
assign g16068 = (g6310&g11775);
assign II31466 = ((~g23821));
assign g8846 = ((~g4779));
assign g9786 = ((~II16832));
assign g5547 = ((~g101));
assign g23385 = ((~g17393)&(~g22517));
assign II18010 = ((~g6369));
assign g21777 = ((~g20228))|((~g6783));
assign g5087 = ((~g1973));
assign g13109 = ((~g9968))|((~g7488));
assign II32958 = ((~g24594));
assign g24869 = (g24047&g18894);
assign II16608 = ((~g5556));
assign g26963 = (g6216&g26539);
assign g15105 = (g4224&g13168);
assign II31068 = ((~g22167));
assign g18521 = ((~g14044));
assign II33358 = ((~g25028));
assign g15531 = ((~II21790));
assign g27258 = ((~g26977)&(~g26257));
assign g28012 = ((~II36513));
assign g16470 = ((~II22512));
assign g25330 = ((~g24873));
assign II27104 = ((~g19239));
assign g25290 = (g24668&g8771);
assign g22773 = ((~II29533));
assign II18752 = ((~g8828));
assign II15818 = ((~g5596));
assign g15819 = ((~g13286))|((~g12392));
assign g11960 = ((~g11252));
assign II23954 = ((~g16154));
assign g13954 = ((~II21012));
assign g7531 = ((~g1180));
assign g25337 = (g24664&g18003);
assign g22873 = ((~II29675));
assign g16974 = ((~g13589));
assign II18172 = ((~g3722));
assign g10624 = (g7195&g5252);
assign g8788 = ((~II15986));
assign g16237 = (g5379&g11886);
assign g30718 = ((~II40444));
assign II32470 = ((~g24058))|((~II32468));
assign g19240 = (g17083)|(g17050)|(II25495);
assign II16241 = ((~g5556));
assign g11630 = ((~g9066)&(~g9081)&(~g9097));
assign g12080 = ((~g10285)&(~g10363)&(~g10430));
assign g5346 = ((~g3106));
assign g24814 = ((~g24239))|((~g24244));
assign g25034 = ((~g23955))|((~g6945));
assign g23597 = ((~II30695));
assign g4650 = ((~g1122));
assign g13605 = ((~g11681));
assign g4321 = ((~II13417));
assign g8681 = ((~II15879));
assign g13073 = ((~g10793));
assign II30841 = ((~g22101));
assign II36732 = ((~g27567))|((~II36731));
assign g23217 = ((~II30104));
assign II29107 = ((~g21435));
assign II23739 = ((~g13548));
assign g27092 = (g5153&g26434);
assign g30684 = ((~g16455)&(~g30337));
assign g8557 = (g3722&g2339);
assign II24092 = ((~g13886))|((~II24091));
assign g21259 = (g20299&g16722&g16682);
assign g30840 = ((~II40772));
assign g21956 = ((~II28494));
assign II23785 = ((~g13551));
assign II39252 = ((~g29695));
assign g4179 = ((~g2106));
assign g15771 = ((~II22019));
assign g30366 = ((~II39909));
assign g20617 = ((~II27176));
assign g5217 = ((~g2673));
assign II31646 = ((~g23692));
assign g13861 = ((~g11613));
assign g18129 = (g5190&g15685);
assign g27780 = ((~II36217));
assign II30663 = ((~g22044));
assign g4601 = ((~g444));
assign g6200 = ((~g542));
assign g27009 = (g23368&g26582);
assign g26629 = ((~g25741));
assign g16639 = (g15210&g15274);
assign II40654 = ((~g30573));
assign g10594 = (g3806&g2667);
assign gbuf30 = (g454);
assign g30103 = (g29869&g11358);
assign II14874 = ((~g1309));
assign II17122 = ((~g7195));
assign g26312 = (g25915&g9610);
assign g15848 = ((~g12657))|((~g6574));
assign g20381 = ((~g17496));
assign g27347 = ((~g27108)&(~g26493));
assign g15790 = ((~g13011));
assign g13240 = ((~g9936));
assign II27969 = ((~g19162));
assign g18891 = ((~g15461));
assign g19218 = ((~II25459));
assign g18548 = ((~g14249)&(~g16082));
assign g12103 = ((~g11450));
assign g26183 = ((~g25957)&(~g13270));
assign g27212 = ((~II35473));
assign g16250 = (g519&g11895);
assign II16954 = ((~g3774));
assign g12920 = ((~g8490)&(~g8506)&(~g8521));
assign g26455 = (g5207&g25808);
assign II17097 = ((~g7936));
assign II31658 = ((~g23785));
assign g22942 = ((~g21263))|((~g2151));
assign g27126 = ((~II35313));
assign g24780 = (g9649&g24132);
assign g4221 = ((~g426));
assign II24226 = ((~g6427))|((~g14316));
assign II32979 = ((~g24598));
assign g22278 = ((~g20722));
assign II39856 = ((~g30276));
assign g10581 = (g7195&g5179);
assign g30286 = ((~g16449)&(~g29982));
assign g28850 = (g27875&g28617);
assign II40757 = ((~g30667));
assign g13847 = (g7521&g12646);
assign g24811 = (g9941&g24161);
assign g25137 = ((~II32889));
assign g22766 = ((~II29516));
assign g22133 = ((~II28671));
assign g26211 = ((~II34135));
assign g28722 = (g28523&g16694);
assign II18713 = ((~g8877));
assign g9956 = (g7085&g4194);
assign II36533 = ((~g27277));
assign g23307 = ((~II30374));
assign g10438 = (g3366&g4908);
assign g22292 = (g21726&g12321);
assign II31682 = ((~g24240));
assign g11723 = ((~g9822))|((~g3678));
assign g25835 = ((~g24742)&(~g24536));
assign g19198 = ((~II25429));
assign g26846 = ((~II34997));
assign g5995 = ((~g2200));
assign II17995 = ((~g6232));
assign g30147 = ((~g30013));
assign II21292 = ((~g11888));
assign II38401 = ((~g28725));
assign II30854 = ((~g22104));
assign g29293 = ((~II38428));
assign g7157 = ((~g453));
assign II20691 = ((~g13327));
assign g30618 = ((~g30412)&(~g25449));
assign g8550 = ((~g3554))|((~g3522));
assign g14067 = (g7703&g12940);
assign g14413 = ((~g12114));
assign II30089 = ((~g22677));
assign II36316 = ((~g15952))|((~II36314));
assign g20190 = (g18415&g9227);
assign g10748 = (g7488&g5385);
assign g30738 = ((~II40498));
assign g14259 = ((~II21137));
assign II37200 = ((~g27907));
assign II17662 = ((~g6425));
assign g22219 = ((~II28781));
assign g14765 = ((~II21301));
assign II40943 = ((~g30834));
assign g25181 = (g24636&g20673);
assign g14359 = ((~g12083));
assign II35715 = ((~g26859))|((~II35714));
assign g26319 = (g4740&g25576);
assign II15949 = ((~g7053));
assign g30528 = ((~II40164));
assign g23631 = (g4168&g22530);
assign g21883 = ((~g19890));
assign g22552 = ((~II29110));
assign g22103 = ((~g21363)&(~g19656));
assign g23796 = (g22739&g17767);
assign g23793 = ((~II31011));
assign g8978 = ((~II16292));
assign g5330 = ((~g1424));
assign g30574 = ((~g30400));
assign g22244 = (g21742&g12198);
assign g16400 = (g1900&g12058);
assign g12215 = ((~g10459)&(~g10521)&(~g10583));
assign g20879 = ((~g19601)&(~g17396));
assign g30006 = (g29928&g22310);
assign g29498 = ((~II38811))|((~II38812));
assign g15740 = (g5319&g13304);
assign g22214 = (g21907&g12045);
assign g23261 = ((~II30236));
assign g28643 = ((~g27942));
assign II19869 = ((~g8726));
assign g25975 = (g24606&g21917);
assign g28578 = ((~g26039)&(~g27734));
assign g23674 = (g22915&g20413);
assign g27792 = ((~II36237));
assign g21821 = (g18753)|(g20309)|(g20294)|(g18668);
assign g18329 = (g5320&g15771);
assign g24225 = ((~g17021)&(~g22281));
assign g28755 = ((~II37716));
assign II27411 = ((~g19457));
assign g25546 = ((~II33374));
assign g25952 = ((~g24735));
assign g15031 = (g4111&g13159);
assign g22209 = ((~II28766))|((~II28767));
assign g10999 = ((~II17904));
assign II26980 = ((~g17086));
assign g21407 = ((~g20499)&(~g13316));
assign II29817 = ((~g21470));
assign g24630 = ((~II32210));
assign g23203 = ((~II30062));
assign g21884 = ((~g19260)&(~g19284));
assign g24887 = ((~II32608))|((~II32609));
assign g27243 = ((~g26802)&(~g10340));
assign g13982 = ((~g11874));
assign g26379 = (g4945&g25669);
assign g11694 = ((~g9968))|((~g3834));
assign g18757 = ((~g14963));
assign g22001 = ((~g21270)&(~g21283));
assign II27321 = ((~g19335));
assign g28418 = ((~g24723)&(~g27846));
assign g26230 = ((~II34168));
assign g13375 = ((~g11481)&(~g11332)&(~g7928)&(~g7880));
assign g24794 = (g2746&g24146);
assign g5234 = ((~II13820));
assign g8167 = ((~II15392));
assign II39349 = ((~g29728))|((~II39347));
assign g28087 = (g27613&g10161);
assign g27868 = ((~g23742)&(~g27632));
assign II24426 = ((~g7134))|((~g14332));
assign II39454 = ((~g29940));
assign g5924 = ((~II14384));
assign g26130 = ((~g23748))|((~g25386));
assign II37319 = ((~g28149));
assign g13267 = ((~II20320));
assign g30806 = ((~II40670));
assign g21561 = ((~II28093));
assign II30516 = ((~g23058));
assign II34872 = ((~g26217));
assign g25081 = ((~g23423)&(~g22202));
assign g9351 = ((~II16566));
assign II22886 = ((~g15661))|((~II22884));
assign g22540 = ((~II29090));
assign g24465 = ((~g23748))|((~g3618));
assign g7156 = ((~g461));
assign g30821 = ((~II40715));
assign g23600 = (g4044&g22490);
assign g22140 = ((~g21398)&(~g19720));
assign g17340 = ((~g16136)&(~g16183));
assign g16047 = (g12130&g10895);
assign g10524 = (g7230&g5095);
assign g25640 = ((~II33463));
assign g17836 = (g4791&g15480);
assign II28527 = ((~g21407));
assign II25294 = ((~g17124));
assign g26892 = ((~g25699))|((~g26283))|((~g25569))|((~g25631));
assign g18872 = ((~g15399));
assign g6435 = ((~g2707));
assign g11431 = (g6369&g900);
assign g7487 = ((~II15012));
assign g23607 = ((~II30713));
assign II28038 = ((~g19957));
assign II26615 = (g14797&g18692&g13657);
assign g16287 = ((~g12962));
assign g27977 = ((~II36450));
assign g29504 = ((~II38838));
assign g25482 = (g24480&g17567);
assign g16052 = (g5591&g11765);
assign g22746 = ((~II29472));
assign g9468 = ((~II16644));
assign g10727 = (g7358&g5372);
assign g20350 = ((~g17410));
assign II24346 = ((~g15873));
assign II29493 = ((~g21010));
assign II38190 = ((~g29093));
assign II32445 = ((~g24054))|((~II32443));
assign g22398 = (g2156&g21222);
assign g18277 = ((~II24279))|((~II24280));
assign g19756 = (g4424&g17624);
assign g28119 = ((~II36786));
assign II24656 = ((~g6190))|((~II24655));
assign II32575 = ((~g18155))|((~g24089));
assign g23339 = ((~g22181)&(~g10238));
assign g29364 = ((~g28894));
assign g21133 = ((~g20108)&(~g20132)&(~g20156));
assign g18226 = ((~g14222));
assign g28451 = (g28133&g9320);
assign g22989 = ((~g21415));
assign II25540 = ((~g92))|((~II25539));
assign II23442 = ((~g13495));
assign g16877 = ((~II22852));
assign g29251 = (g28855&g8856);
assign g28703 = ((~II37656));
assign g13045 = ((~g9534))|((~g6912));
assign g28352 = ((~g15624)&(~g28065));
assign g10287 = (g6486&g596);
assign gbuf15 = (g2845);
assign g28744 = ((~g15030)&(~g28439));
assign g15487 = (g4800&g12825);
assign g17092 = ((~g13530));
assign II30299 = ((~g22694));
assign II31790 = ((~g23459));
assign g15759 = ((~g12565))|((~g6314));
assign g30311 = ((~II39776));
assign g12225 = ((~II19401));
assign II28137 = ((~g20067));
assign g26076 = ((~II33974));
assign g12270 = ((~g10535)&(~g10595)&(~g10640));
assign II23264 = ((~g9857))|((~g14413));
assign g19573 = ((~II26006));
assign g26590 = ((~g25609));
assign g12056 = ((~g10225)&(~g10311)&(~g10388));
assign II17840 = ((~g8107));
assign g17398 = (g4026&g15043);
assign II20386 = ((~g10796));
assign II32886 = ((~g24549));
assign g12162 = ((~g10390)&(~g10452)&(~g10515));
assign II29547 = ((~g21031));
assign g22759 = (g14360&g21619);
assign II35419 = ((~g26828));
assign II19859 = ((~g10617));
assign II32829 = ((~g24059));
assign g4997 = ((~g2433));
assign II36432 = ((~g27585));
assign II28130 = ((~g20025));
assign g15459 = (g4897&g13218);
assign II22983 = ((~g14106))|((~II22981));
assign g10229 = ((~g5349));
assign II35351 = ((~g26272));
assign g20802 = ((~II27391));
assign g19262 = ((~II25540))|((~II25541));
assign g11541 = ((~II18599));
assign g28275 = ((~II37074));
assign II15192 = ((~g2959))|((~II15190));
assign g28153 = ((~g27397));
assign g11871 = ((~g11105));
assign g19676 = (g2072&g18832);
assign g15666 = (g5233&g13268);
assign II23619 = ((~g13535));
assign g24108 = ((~g22434));
assign g26817 = ((~g15375)&(~g26317));
assign g27762 = ((~g27530)&(~g27091));
assign g20700 = ((~g20153))|((~g2903));
assign II18824 = ((~g9084));
assign g17991 = ((~g14450));
assign g19358 = ((~II25768));
assign g20594 = ((~II27107));
assign g5973 = ((~g2321));
assign II36860 = ((~g27386));
assign g26035 = (g25523&g19483);
assign gbuf63 = (g528);
assign g13445 = ((~II20634));
assign g30001 = (g29897&g8449);
assign g19666 = (g1326&g18825);
assign g29321 = (g29008&g28979);
assign g6314 = ((~II14734));
assign g13059 = ((~g9534))|((~g6912));
assign II24710 = ((~g14502))|((~II24709));
assign g26171 = (g2059&g25942);
assign g22721 = ((~g21164));
assign g24429 = (g24115&g13614);
assign g6368 = ((~II14739));
assign g13344 = ((~II20421));
assign II26469 = ((~g16672));
assign g27321 = ((~g27063)&(~g26416));
assign g9092 = (g6448&g7673);
assign g17065 = (g3566&g10735&g14381);
assign g30542 = ((~II40206));
assign II25272 = ((~g17051));
assign II20339 = ((~g9084));
assign g23843 = (g22966&g9734);
assign g28483 = ((~g27776));
assign g20352 = ((~g17416));
assign II15942 = ((~g6945));
assign g11621 = ((~II18800))|((~II18801));
assign g20948 = ((~g19735)&(~g15336));
assign g8327 = (g3254&g219);
assign gbuf167 = (g2003);
assign g4067 = ((~g1555));
assign II28473 = ((~g21030));
assign g23667 = (g22644&g20408);
assign g16625 = (g15118&g15188);
assign II24111 = ((~g13963))|((~II24110));
assign g19672 = (g4162&g17471);
assign g30486 = (g30171&g11376);
assign g9202 = ((~II16482));
assign g26544 = ((~g25479));
assign g13631 = (g6189&g12481);
assign g12318 = ((~II19485));
assign g14420 = ((~II21190));
assign g28807 = ((~II37768));
assign g11102 = ((~II18016));
assign g20534 = ((~g18505));
assign g10308 = (g3566&g4674);
assign g11522 = ((~II18542));
assign g22470 = ((~II29016));
assign g27057 = (g23377&g26623);
assign g29583 = ((~II38975));
assign g15681 = (g5256&g13279);
assign g27986 = ((~II36459));
assign g29408 = ((~II38609));
assign g9488 = ((~g5914));
assign g23818 = (g22900&g17788);
assign II24603 = ((~g14135))|((~II24601));
assign g13152 = ((~g9196));
assign g24870 = (g18281&g23786);
assign g27589 = ((~g27168));
assign g3650 = ((~II13211));
assign II33488 = ((~g25054));
assign gbuf5 = (g2870);
assign g29618 = ((~g13997)&(~g29261));
assign g5003 = ((~g2510));
assign II32126 = ((~g24212));
assign II30979 = ((~g22143));
assign II33667 = ((~g24470));
assign II16218 = ((~g5473));
assign g26247 = ((~II34195));
assign g14747 = ((~g12324));
assign g16347 = (g5900&g11982);
assign g10447 = (g7162&g4933);
assign II15989 = ((~g6053));
assign g11910 = ((~g11166));
assign II28461 = ((~g20998));
assign g21925 = (g19384&g11749);
assign g19267 = (g16924&g14395&g14301);
assign II22563 = ((~g14830));
assign II30104 = ((~g22760));
assign g28740 = ((~g28488));
assign g24879 = ((~II32583));
assign g9776 = (g3410&g4029);
assign gbuf204 = (g2646);
assign g6167 = ((~g2052));
assign II37590 = ((~g28555));
assign g22366 = ((~g20827));
assign g25277 = (g24648&g8714);
assign g4095 = ((~g130));
assign g14830 = ((~II21329));
assign g22431 = ((~II28975));
assign g15436 = (g4868&g13213);
assign g26137 = ((~g6068)&(~g24183)&(~g25355));
assign g27260 = ((~g26979)&(~g26259));
assign g30459 = ((~II40021));
assign g27883 = ((~g6087)&(~g27632)&(~g25361));
assign gbuf116 = (g1244);
assign g29754 = ((~g16178)&(~g29607));
assign g20775 = ((~g20228))|((~g3566));
assign II30389 = ((~g22225));
assign g10301 = (g6751&g4652);
assign g27141 = ((~g26251));
assign g4240 = ((~g849));
assign g15580 = (g5121&g13242);
assign g27004 = (g23344&g26574);
assign g27689 = ((~II36078));
assign g24544 = ((~II32074));
assign g30509 = ((~II40107));
assign II15245 = ((~g2941))|((~II15244));
assign g23201 = ((~II30056));
assign II18369 = ((~g4325))|((~II18368));
assign g25300 = (g24687&g8794);
assign g30741 = ((~II40507));
assign g11438 = ((~II18402));
assign g28606 = ((~g26040)&(~g27737));
assign II14246 = ((~g3227));
assign II41053 = ((~g30939));
assign II33491 = ((~g24501));
assign II26931 = ((~g17340));
assign II23093 = ((~g9326))|((~g13935));
assign g19557 = (g8053&g17249);
assign g14023 = (g7682&g12922);
assign g10730 = ((~g6173));
assign g13063 = ((~g10835));
assign g26574 = ((~g25562));
assign g12988 = ((~II20032))|((~II20033));
assign g19888 = (g18247&g16180);
assign g11700 = ((~g9968))|((~g3834));
assign g16654 = ((~g14690)&(~g12477));
assign II40527 = ((~g30691));
assign II36718 = ((~g27327));
assign g21426 = ((~II27969));
assign g26254 = ((~II34210));
assign g5053 = ((~g1271));
assign g17695 = (g4549&g15357);
assign g5854 = ((~g252));
assign g26580 = ((~g25579));
assign g5847 = (g2400&g2454);
assign g12097 = ((~g10301)&(~g10377)&(~g10441));
assign g24838 = (g12945&g24175);
assign g17618 = (g4412&g15287);
assign II29235 = ((~g20918));
assign g24860 = ((~II32519))|((~II32520));
assign II33514 = ((~g25039));
assign g6838 = ((~II14842));
assign g9449 = ((~II16630));
assign g29084 = ((~II38053));
assign II27667 = ((~g20507));
assign g24775 = (g15694&g24128);
assign g21373 = (g9488&g20372);
assign g12940 = ((~g8980));
assign g18949 = ((~g15685));
assign g15471 = ((~II21730));
assign g20506 = (g17499&g12025);
assign II38761 = ((~g29281));
assign II20455 = ((~g8578));
assign g18860 = ((~g15360));
assign g13177 = ((~g9371));
assign g20347 = ((~g17399));
assign g16939 = (g7158&g15129);
assign II34701 = ((~g26193));
assign g23083 = ((~g21160)&(~g21193));
assign II25071 = ((~g14910));
assign g13671 = (g6418&g12521);
assign g6162 = ((~g1240));
assign g15594 = (g5148&g13249);
assign II16703 = ((~g6751));
assign g29053 = ((~g9264))|((~g28567));
assign g3252 = ((~II13152));
assign g8375 = ((~II15577));
assign II26444 = ((~g17076));
assign II33723 = ((~g24477));
assign g15832 = ((~g12565))|((~g6232));
assign g13927 = ((~g12789));
assign II18362 = ((~g5837));
assign g22405 = ((~II28949));
assign g25319 = ((~g24857));
assign g11893 = ((~g11138));
assign II19657 = ((~g10839));
assign II22852 = ((~g13600));
assign g24982 = ((~g23505));
assign g14796 = ((~II21321));
assign II36900 = ((~g28023));
assign g17303 = ((~g16105)&(~g16137));
assign g24790 = (g9795&g24142);
assign g15335 = (g4489&g12749);
assign g4545 = ((~g1807));
assign II24732 = ((~g13633));
assign g20163 = ((~g17973));
assign II31649 = ((~g23738));
assign II18133 = ((~g6448));
assign II20264 = ((~g9027));
assign g27221 = ((~II35500));
assign II32480 = ((~g24065))|((~II32478));
assign II35452 = ((~g27161));
assign g28371 = ((~g15793)&(~g28127));
assign g5424 = ((~II13984));
assign II33655 = ((~g24527));
assign g29334 = ((~II38515));
assign II37906 = ((~g28556));
assign g13839 = (g7557&g12643);
assign II18256 = ((~g6574));
assign g30396 = (g30237&g9013);
assign g23185 = ((~II30008));
assign g4606 = ((~g579));
assign g23585 = ((~II30669));
assign g25207 = ((~g24747)&(~g23551));
assign g26029 = (g25445&g24952);
assign g11274 = ((~II18220));
assign II35536 = ((~g26844));
assign g28642 = ((~g27939));
assign g24540 = (g18548&g23089&g23403);
assign g12038 = ((~g11361));
assign g29531 = (g29202&g29371);
assign g29520 = (g28731&g29361);
assign g19108 = (g18744&g15003&g16371&g13825);
assign II21282 = ((~g11675));
assign g30378 = ((~II39939));
assign g18862 = ((~g15376));
assign II34857 = ((~g26355));
assign g10472 = (g7391&g2645);
assign g28443 = ((~II37394));
assign g30581 = ((~II40297));
assign g3773 = ((~g2380));
assign g29998 = (g29922&g22278);
assign g14053 = ((~g12866));
assign g4332 = ((~g134));
assign II14731 = ((~g135));
assign II25922 = ((~g2151))|((~II25921));
assign g19939 = (g16583&g16954&g16560);
assign II25740 = ((~g1439))|((~g17842));
assign II20382 = ((~g10907));
assign II22382 = ((~g520));
assign g19291 = ((~II25612));
assign II16209 = ((~g5438));
assign g20970 = ((~g19769)&(~g15403));
assign II38094 = ((~g28363));
assign II16476 = ((~g6448));
assign g29326 = ((~II38499));
assign g6140 = ((~g524));
assign g7928 = ((~g3204));
assign g15995 = ((~g12926))|((~g6980));
assign g19901 = (g1372&g18947);
assign II26458 = ((~g17985));
assign II32355 = ((~g18014))|((~g24003));
assign g22282 = (g21752&g12299);
assign g19604 = (g3948&g17354);
assign g12378 = ((~g10847));
assign II40266 = ((~g30365));
assign g16072 = (g12275&g10924);
assign g24332 = ((~II31670));
assign II20559 = ((~g11937));
assign g5987 = ((~II14459));
assign g22600 = ((~II29180));
assign II40589 = ((~g30622))|((~II40587));
assign g23709 = (g22826&g17591);
assign II37357 = ((~g27824))|((~II37356));
assign g6157 = ((~g686));
assign II29481 = ((~g21007));
assign II36132 = ((~g27366));
assign II37581 = ((~g28374));
assign g23954 = ((~g4632)&(~g22987));
assign g27827 = ((~g6087)&(~g27632)&(~g25314));
assign g6294 = ((~g1937));
assign II29132 = ((~g21781));
assign g10493 = (g6643&g5030);
assign II30407 = ((~g22970));
assign II30944 = ((~g22132));
assign g26275 = ((~g25315));
assign g3805 = ((~g2384));
assign g16984 = (g7538&g15236);
assign g29355 = ((~g29128)&(~g17065));
assign g15534 = ((~II21793));
assign g24072 = ((~g22004)&(~g20826));
assign g23219 = ((~II30110));
assign II28360 = ((~g20163));
assign g22088 = ((~g21350)&(~g19631));
assign g17138 = (g7676&g14068);
assign g16998 = (g7862&g15353);
assign g24495 = ((~g23717)&(~g19783));
assign II13916 = ((~g1033));
assign g11268 = ((~II18214));
assign g11963 = ((~g11259));
assign g11039 = ((~II17954));
assign g23236 = ((~II30161));
assign g11909 = ((~g11163));
assign g15591 = (g5018&g12868);
assign II38074 = ((~g28356));
assign II24271 = ((~g6180))|((~g13922));
assign g23295 = ((~II30338));
assign II32568 = ((~g18131))|((~II32567));
assign g29091 = ((~II38068));
assign g27483 = ((~II35829));
assign g21068 = (g20058&g14194&g14280);
assign g13167 = ((~g9303));
assign g22483 = (g646&g21861);
assign g25694 = ((~II33520));
assign g20271 = (g18679&g14910&g16351);
assign g29244 = ((~II38339));
assign g14132 = ((~g8911))|((~g12527))|((~g12515));
assign II27408 = ((~g19431));
assign g4786 = ((~g1276));
assign g23561 = ((~II30623));
assign g29153 = ((~II38202));
assign g13903 = ((~g11815));
assign II33548 = ((~g25064));
assign g27565 = ((~g26768)&(~g19100));
assign g25234 = ((~g24789)&(~g23605));
assign II20465 = ((~g11330))|((~g11263));
assign II33680 = ((~g24471));
assign g12699 = ((~II19791));
assign g20883 = ((~g19615)&(~g17409));
assign II20283 = ((~g9050));
assign II20544 = ((~g11628));
assign II24319 = ((~g14217))|((~II24317));
assign g22199 = (g16164)|(g20858);
assign g21026 = ((~g19861)&(~g17966));
assign g16343 = (g5895&g11969);
assign II40949 = ((~g30835));
assign g25104 = ((~g23832));
assign g30098 = (g29853&g11284);
assign g27044 = (g22016&g26610);
assign g24043 = ((~g23033)&(~g7455));
assign g18568 = ((~II24656))|((~II24657));
assign g25012 = ((~g23644))|((~g6448));
assign g27296 = ((~g27030)&(~g26363));
assign g11875 = ((~g9811)&(~g9926)&(~g10062));
assign g27338 = ((~g27090)&(~g26457));
assign g20806 = ((~II27395));
assign g8533 = ((~g3398))|((~g3366));
assign g9584 = (g6369&g8221);
assign g6298 = ((~g2013));
assign g9916 = ((~II16918));
assign g14322 = ((~g12959));
assign g28654 = ((~g27770)&(~g27355));
assign II25966 = ((~g16654));
assign g27731 = (g27470&g19383);
assign g15219 = (g4405&g13181);
assign g30300 = ((~g13502)&(~g30001));
assign II24352 = ((~g14238))|((~II24351));
assign g16797 = ((~g15080));
assign II38068 = ((~g28354));
assign g8676 = (g6643&g7838);
assign II36927 = ((~g28048));
assign g19025 = ((~II25138));
assign g12886 = (g9534)|(g3398);
assign g28342 = ((~g15460)&(~g28008));
assign g15913 = ((~g11647));
assign g20193 = ((~g18691));
assign g7535 = ((~g2555));
assign g17802 = ((~g13907));
assign g14263 = ((~g12941));
assign g27182 = (g26151&g22217);
assign g28529 = (g27743)|(g25818);
assign II14593 = ((~g1765));
assign g26803 = ((~g15105)&(~g26213));
assign g26755 = (g26083&g22239);
assign g12124 = ((~g10353)&(~g10413)&(~g10475));
assign II25940 = ((~g18142))|((~II25938));
assign g11600 = ((~g9049)&(~g9064)&(~g9078));
assign g30032 = ((~g24712)&(~g29927));
assign g4967 = ((~g2095));
assign g30331 = ((~II39832));
assign II14891 = ((~g1925));
assign II26115 = ((~g16845));
assign II41108 = ((~g30967));
assign g30226 = (g30048&g9041);
assign g30748 = ((~II40524));
assign g17025 = ((~g15904)&(~g15880)&(~g15859));
assign g19104 = (g13687&g16302&II25291);
assign II17059 = ((~g6637))|((~g6309));
assign g24360 = ((~II31754));
assign g28313 = ((~II37188));
assign II16047 = ((~g6063));
assign g21590 = ((~II28119));
assign g9727 = ((~II16776));
assign g22901 = ((~II29694));
assign g20249 = (g18679&g18758&g13687&g16351);
assign g26047 = ((~g25619)&(~g24902));
assign II32451 = ((~g18038))|((~g24056));
assign g15871 = ((~g12711))|((~g6838));
assign g10402 = (g7085&g4854);
assign g12120 = ((~g10327)&(~g10404)&(~g10467));
assign g16802 = ((~g13469)&(~g3897));
assign II33297 = ((~g24430));
assign g11263 = ((~II18198))|((~II18199));
assign g16856 = (g6443&g14794);
assign g26490 = ((~II34456));
assign II23824 = ((~g14904));
assign II31538 = ((~g23775));
assign g29579 = ((~g29399)&(~g17001));
assign II27785 = ((~g20064));
assign II33714 = ((~g24547));
assign II32546 = ((~g17903))|((~g23906));
assign II15230 = ((~g499));
assign II17878 = ((~g8031));
assign g29113 = ((~g28381)&(~g8907));
assign g19316 = (g18063&g3110);
assign g9364 = (g3254&g8053);
assign g9013 = ((~II16335));
assign g9633 = (g3254&g3931);
assign g26834 = ((~II34971));
assign g30493 = ((~II40075));
assign g21951 = ((~II28479));
assign g20460 = (g17351&g13644);
assign II34461 = ((~g25280));
assign II24703 = ((~g7259))|((~II24702));
assign g13330 = ((~g10357));
assign g12043 = ((~g10210)&(~g10296)&(~g10372));
assign g30795 = ((~II40643));
assign g14381 = ((~II21178));
assign II34842 = ((~g26505));
assign II28997 = ((~g21759));
assign g10570 = (g3522&g5164);
assign g4933 = ((~g1404));
assign g25377 = (g24700&g18324);
assign g20091 = (g16804&g3136);
assign g27189 = ((~II35404));
assign g18023 = (g5067&g15615);
assign g27906 = ((~g16127)&(~g27656));
assign gbuf144 = (g1768);
assign g17159 = ((~g14642))|((~g14657));
assign g20983 = ((~g19797)&(~g17797));
assign g26874 = ((~II35058))|((~II35059));
assign g16218 = (g5777&g11877);
assign g28771 = ((~g15218)&(~g28463));
assign g27521 = ((~g26766)&(~g24439));
assign g25280 = ((~g24924)&(~g18164));
assign II39460 = ((~g29932));
assign g15247 = (g4479&g13187);
assign g26795 = ((~g26050)&(~g10340));
assign II40125 = ((~g30466));
assign g7754 = ((~g322));
assign II29539 = ((~g21028));
assign g25561 = (g24495&g20462);
assign g23589 = ((~II30679));
assign II40176 = ((~g30331));
assign II25189 = ((~g19008));
assign g30909 = ((~II40979));
assign g28972 = ((~II37939));
assign II34392 = ((~g25266));
assign g22248 = ((~g20662));
assign g25725 = ((~g24731)&(~g24512));
assign g28038 = ((~II36571));
assign g16722 = ((~g14895));
assign g28408 = (g7806&g27861);
assign II20886 = ((~g12499));
assign g29360 = ((~g28871));
assign g28843 = (g27834&g28581);
assign g17278 = ((~II23364));
assign g4162 = ((~g1539));
assign II20430 = ((~g11262))|((~II20429));
assign g12235 = ((~g8294));
assign g23057 = ((~g21599));
assign g29926 = ((~g29718)&(~g22367));
assign g25138 = ((~II32892));
assign g12560 = ((~g8745));
assign II39002 = ((~g29506));
assign g20472 = (g17314&g13669);
assign g7848 = ((~g1890));
assign II36918 = ((~g28025));
assign g26711 = ((~II34740));
assign g10058 = (g3522&g4263);
assign g8643 = ((~II15833));
assign g29396 = ((~g29057));
assign g21456 = (g15296&g20437);
assign II16193 = ((~g5417));
assign II13922 = ((~g1724));
assign g30505 = ((~g14229)&(~g30224));
assign g19716 = (g2033&g18846);
assign II30338 = ((~g22837));
assign g24438 = ((~g23408)&(~g10340));
assign II31928 = ((~g24255));
assign g5915 = ((~g2303));
assign II15571 = ((~g7085));
assign g17679 = ((~II23763));
assign II29333 = ((~g20953));
assign g16030 = (g7667&g11746);
assign g27612 = ((~g27184)&(~g17065));
assign g9309 = ((~II16544));
assign g21448 = (g15210&g20431);
assign g17631 = (g6435&g15308);
assign g17409 = (g4052&g15052);
assign g21137 = (g5750&g19272);
assign g28054 = ((~II36615));
assign g5609 = ((~g1201));
assign g21159 = (g19524)|(g16578)|(g14301);
assign g23278 = ((~II30287));
assign g11686 = ((~g9822))|((~g3678));
assign g23558 = (g8200&g22422);
assign II38104 = ((~g28367));
assign g19886 = (g2740&g18940);
assign g11462 = ((~II18426));
assign g5246 = ((~g1830));
assign g30012 = ((~g29523)&(~g29945));
assign g16181 = ((~II22317))|((~II22318));
assign g28162 = ((~g27432));
assign II25549 = (g17190)|(g17175)|(g17165);
assign II16677 = ((~g3306));
assign g21972 = ((~g20914)&(~g10238));
assign g23243 = ((~II30182));
assign g12962 = ((~II20009));
assign g20858 = ((~g19491));
assign II27585 = ((~g20376));
assign g12339 = ((~g10650)&(~g10678)&(~g10704));
assign g28405 = (g7796&g27847);
assign II29863 = ((~g21346));
assign II21632 = ((~g13093));
assign g10232 = ((~II17206));
assign II40901 = ((~g30725));
assign g5101 = ((~g2116));
assign g20178 = ((~g16842));
assign g22693 = ((~II29351));
assign g29080 = ((~g9407))|((~g28595));
assign g5655 = ((~g813));
assign II27044 = ((~g19247));
assign II15277 = ((~g2935))|((~II15276));
assign g15170 = ((~g12125));
assign II33670 = ((~g25066));
assign II27531 = ((~g20343));
assign g10326 = (g7085&g4714);
assign II16163 = ((~g6031));
assign II15019 = ((~g2830));
assign g8001 = ((~g830));
assign g16019 = (g5507&g11742);
assign g14139 = ((~g11965));
assign g24398 = ((~II31868));
assign g27156 = ((~II35351));
assign g26736 = ((~II34815));
assign g26651 = ((~g25838));
assign g11234 = ((~II18160));
assign g7616 = ((~g313));
assign g10709 = (g7230&g5358);
assign g29848 = ((~g29761));
assign II15246 = ((~g2944))|((~II15244));
assign g25202 = ((~g24566)&(~g22907));
assign g25411 = ((~g24842));
assign g24060 = ((~g23040));
assign gbuf126 = (g1831);
assign II13246 = ((~g2987));
assign II15662 = ((~g3722));
assign II40146 = ((~g30344));
assign g29096 = ((~g9649))|((~g28540));
assign g4372 = ((~g1041));
assign g13038 = ((~g9676))|((~g7162));
assign II27717 = (g19345&g19321&g19304);
assign II17300 = ((~g3806));
assign g6118 = ((~II14637));
assign g19636 = (g1378&g18812);
assign g24739 = ((~g23941)&(~g22835));
assign g26718 = ((~II34761));
assign II20643 = ((~g13296));
assign g25861 = ((~g24657)&(~g24546));
assign II35014 = ((~g26498));
assign g5774 = ((~g1439));
assign II27167 = ((~g20457));
assign g23500 = ((~II30544));
assign II29271 = ((~g20752));
assign g29177 = ((~II38258));
assign II15784 = ((~g6000));
assign g23358 = ((~g22227)&(~g18407));
assign g30831 = ((~II40745));
assign g19723 = (g2707&g18850);
assign g17460 = (g4048&g16012);
assign g16466 = ((~g12017));
assign II33343 = ((~g25024));
assign II32309 = ((~g17903))|((~II32308));
assign g25940 = ((~g24428)&(~g17100));
assign II32116 = ((~g24208));
assign g23552 = (g6136&g22415);
assign g26013 = ((~II33891));
assign g26570 = ((~g25549));
assign II36243 = ((~g27587));
assign g18354 = ((~II24362))|((~II24363));
assign II15932 = ((~g5423));
assign g15346 = ((~II21615));
assign g22260 = ((~g20684));
assign II14860 = ((~g626));
assign g22299 = ((~g21773)&(~g20104));
assign g21724 = ((~g20228))|((~g6783));
assign g22598 = ((~II29174));
assign g23392 = ((~g17460)&(~g22557));
assign g24557 = ((~g15699)&(~g23942));
assign g18201 = ((~g16123)&(~g6568));
assign g28526 = ((~II37471));
assign II27020 = ((~g19182));
assign g23691 = ((~II30857));
assign g24531 = ((~II32057));
assign II32931 = ((~g24872));
assign g19098 = ((~II25283));
assign g13422 = ((~II20565));
assign II40877 = ((~g30812));
assign II20836 = ((~g13182));
assign g16809 = ((~g15842));
assign II32719 = ((~g23359));
assign g23399 = ((~g17506)&(~g22581));
assign g26320 = (g25852)|(g25870);
assign II18381 = ((~g6232));
assign g9806 = (g3566&g4055);
assign II36524 = ((~g27275));
assign g27063 = (g23388&g26629);
assign II13176 = ((~g630));
assign g7745 = ((~g2391));
assign g28718 = (g28473&g19380);
assign g24848 = ((~II32479))|((~II32480));
assign g26828 = ((~II34957));
assign g23538 = (g5944&g22376);
assign g29302 = (g29026&g28928);
assign g23569 = ((~II30639));
assign II25383 = ((~g18755));
assign g19280 = ((~g16596));
assign g15421 = (g4665&g12791);
assign g29785 = ((~g29485)&(~g29238));
assign g11927 = ((~g10987));
assign g24239 = (g19387)|(g22401);
assign g30582 = ((~II40300));
assign II16318 = ((~g5556));
assign g22802 = ((~II29588));
assign g28291 = ((~II37122));
assign g26900 = ((~II35099));
assign II26508 = (g18644&g18637&g18618);
assign II21838 = ((~g11712));
assign g25841 = ((~II33683));
assign g26612 = ((~g25681));
assign g4598 = ((~g398));
assign g11946 = ((~g10057)&(~g10145)&(~g10217));
assign g23210 = ((~II30083));
assign II17143 = ((~g7303));
assign g28975 = ((~II37942));
assign g25720 = ((~II33548));
assign g29619 = (g29247&g11259);
assign II18190 = ((~g7922))|((~g7895));
assign II38035 = ((~g28345));
assign g10045 = (g3410&g4246);
assign g12007 = ((~g11327));
assign g30130 = ((~II39647));
assign II17913 = ((~g7015));
assign g17871 = ((~II23932));
assign g8024 = ((~g2842));
assign g28363 = ((~g15739)&(~g28111));
assign g16940 = ((~II22893));
assign g21589 = (g3002&g19890);
assign II17637 = ((~g6204));
assign g11290 = ((~II18238));
assign g23901 = ((~II31171));
assign II18305 = ((~g6314));
assign II36663 = ((~g27313));
assign g24550 = (g18548&g23420&g19948);
assign II18435 = ((~g5635));
assign II39691 = ((~g30034))|((~II39689));
assign g26262 = (g25899&g9446);
assign II18500 = ((~g8924));
assign g11807 = ((~g9584)&(~g9664)&(~g9779));
assign II16328 = ((~g3900));
assign g29376 = ((~g28959));
assign g9748 = (g6838&g3990);
assign g24598 = ((~II32178));
assign g18859 = ((~g15357));
assign II30626 = ((~g22034));
assign g11105 = ((~II18019));
assign g16263 = (g5821&g11908);
assign g11414 = ((~II18378));
assign g29857 = ((~g29676));
assign II39059 = ((~g29561));
assign g6057 = ((~II14550));
assign g23623 = (g4139&g22523);
assign g26634 = ((~g25755));
assign II36639 = ((~g27306));
assign g27774 = (g5702&g27361);
assign g6447 = ((~II14760));
assign g23731 = ((~II30917));
assign g25266 = ((~g24881)&(~g17912));
assign g8511 = (g3722&g2312);
assign g10212 = (g5473&g1125);
assign g28147 = ((~g27655)&(~g17065));
assign II33249 = ((~g24890));
assign g16379 = (g2592&g12007);
assign g6486 = ((~II14769));
assign g28222 = ((~II36915));
assign II39255 = ((~g29698));
assign g29955 = (g29787&g28993);
assign g16482 = ((~II22548));
assign g11743 = ((~g8530));
assign II22536 = ((~g14829));
assign g26579 = ((~g25576));
assign g16506 = ((~II22599));
assign g4471 = ((~g384));
assign g23134 = ((~II29881));
assign g10115 = (g6678&g4357);
assign g10937 = ((~II17834));
assign II33621 = ((~g24465));
assign g27172 = ((~g26485));
assign g20976 = ((~g19778)&(~g15422));
assign g17214 = ((~g13585));
assign g25355 = ((~g24797));
assign g25461 = (g6190&g24805);
assign II29606 = ((~g21364));
assign g24288 = ((~II31538));
assign g12294 = ((~g8475));
assign II18470 = ((~g8808));
assign II19894 = ((~g10744));
assign II33335 = ((~g25010));
assign g8333 = ((~II15535));
assign g24872 = ((~II32556));
assign II27188 = ((~g20441));
assign g25519 = ((~II33347));
assign g27319 = ((~g27061)&(~g26414));
assign g9927 = (g6574&g4171);
assign g10834 = ((~II17681));
assign II24454 = ((~g14450))|((~II24452));
assign g28303 = ((~II37158));
assign II35527 = ((~g26900));
assign g27219 = ((~II35494));
assign g17098 = ((~g14747));
assign II15657 = ((~g6838));
assign g19788 = (g4558&g17698);
assign g27710 = ((~II36141));
assign g22334 = ((~g20799));
assign g8295 = ((~g3617));
assign g23861 = ((~II31109));
assign g28175 = ((~g27498));
assign g29835 = ((~g29667));
assign II37928 = ((~g28556));
assign g19228 = (g16662&g12125);
assign g19746 = (g4392&g17604);
assign g14097 = (g7706&g12943);
assign II33136 = ((~g24986));
assign g13228 = ((~g8841)&(~g8861)&(~g8892));
assign II14976 = ((~g2006));
assign II32678 = ((~g23823))|((~II32677));
assign II32506 = ((~g23324));
assign II34479 = ((~g25202));
assign g16608 = ((~II22657));
assign g15366 = ((~g11917));
assign II27038 = ((~g20082));
assign g5813 = ((~g921));
assign g12503 = ((~g8278))|((~g5438));
assign g10930 = ((~II17813));
assign g27577 = ((~g4985)&(~g26901));
assign II15856 = ((~g3522));
assign g19188 = (g17830)|(g18096);
assign g20340 = ((~g17372));
assign g19841 = (g686&g18911);
assign g7957 = ((~g481));
assign g13161 = ((~g9257));
assign g30191 = ((~g30024));
assign g5594 = ((~g793));
assign g30714 = ((~II40432));
assign II18350 = ((~g7195));
assign g27525 = ((~II35897));
assign II16128 = ((~g6103));
assign II34363 = ((~g25930));
assign g19116 = (g13774&g16404&II25311);
assign g16088 = ((~g12816));
assign g24511 = ((~g15411)&(~g23831));
assign II14675 = ((~g1905));
assign g16101 = (g6197&g11794);
assign II17984 = ((~g7976));
assign g26066 = ((~g25431))|((~g25395))|((~g25283));
assign g10651 = (g3494&g1306);
assign g30984 = ((~II41126));
assign II27297 = ((~g19390));
assign II40611 = ((~g30708));
assign g23283 = ((~II30302));
assign g15618 = ((~g9391))|((~g9216))|((~g12857));
assign g30983 = ((~II41123));
assign g14374 = ((~g12099));
assign II31697 = ((~g23791));
assign g22678 = ((~II29326));
assign g8662 = ((~II15856));
assign II34210 = ((~g25761));
assign g19203 = (g18290)|(g18363);
assign II34108 = ((~g25222));
assign g30609 = ((~g30412)&(~g2606));
assign g5738 = ((~II14182));
assign II30800 = ((~g22088));
assign g12830 = ((~II19891));
assign g10967 = ((~II17860));
assign g24178 = ((~g16908)&(~g22211));
assign II17892 = ((~g6232));
assign g12743 = ((~g8817));
assign g30965 = ((~g30959));
assign g17375 = ((~II23463));
assign II39074 = ((~g29556));
assign II40560 = ((~g30597))|((~II40558));
assign II39922 = ((~g30295));
assign g16785 = ((~II22768));
assign g20518 = ((~g18466));
assign gbuf137 = (g1733);
assign g19651 = (g4079&g17425);
assign II21361 = ((~g13026));
assign g23800 = ((~II31024));
assign g19522 = (g16913)|(g16728)|(g16686);
assign g14320 = ((~g12061));
assign g21803 = (g19135)|(g16943)|(g14863);
assign g21229 = (g19578&g14797&g16665);
assign g30902 = ((~II40958));
assign g26074 = (g25948&g21144);
assign g23212 = ((~II30089));
assign II18569 = ((~g8867));
assign g10646 = ((~II17557));
assign g19353 = ((~g16651));
assign g30665 = ((~g16368)&(~g30475));
assign g30838 = ((~II40766));
assign g29255 = (g28855&g8885);
assign g8233 = ((~g1551));
assign g27673 = (g26854&g11312);
assign g20110 = (g18070&g9286);
assign g26700 = ((~II34707));
assign g21066 = ((~g20519));
assign g21034 = ((~g19873)&(~g18012));
assign g23915 = (g22980&g10090);
assign g14229 = (g7748&g12980);
assign g21703 = ((~g16629)&(~g20067));
assign g25539 = ((~g25088)&(~g6157));
assign II16990 = ((~g3338));
assign g30880 = ((~II40892));
assign g3236 = ((~II13104));
assign II25240 = ((~g16934));
assign II22706 = ((~g13348))|((~II22705));
assign II28972 = ((~g21736));
assign g28950 = ((~II37917));
assign g30264 = ((~g16348)&(~g30098));
assign g29945 = (g29773&g28894);
assign g25629 = (g3024&g25116);
assign g26637 = ((~g25773));
assign g20481 = ((~g18201))|((~g1332));
assign II29283 = ((~g20937));
assign g26208 = ((~II34128));
assign g13024 = ((~g11481)&(~g8045)&(~g7928)&(~g7880));
assign g9320 = ((~II16549));
assign g15762 = ((~g13011));
assign II19929 = ((~g10728));
assign II18154 = ((~g6945));
assign g27437 = ((~II35777));
assign II34773 = ((~g26247));
assign g10272 = (g3834&g4587);
assign II30164 = ((~g22655));
assign g27613 = ((~g27165));
assign II24298 = ((~g6209))|((~g14028));
assign g20309 = (g15003&g18796&g13774&g16404);
assign g19863 = (g18155&g16130);
assign g20387 = ((~g17520));
assign II27311 = ((~g19401));
assign g28383 = (g740&g27780);
assign g5434 = ((~g3084));
assign g15307 = ((~g12228));
assign g23725 = ((~II30901));
assign g10167 = (g3678&g4418);
assign g14329 = ((~II21160));
assign g25576 = ((~II33399));
assign g10090 = ((~II17054));
assign g30660 = ((~g16324)&(~g30465));
assign II14020 = ((~g1657));
assign g20446 = ((~g17761));
assign g21737 = ((~g20164))|((~g6314));
assign g24603 = (g23518&g23505);
assign g22671 = ((~II29307));
assign g30552 = ((~II40236));
assign g22238 = (g21939&g12181);
assign g13410 = ((~II20529));
assign g26408 = (g5072&g25729);
assign g21104 = ((~g20050)&(~g20085)&(~g20106));
assign g20813 = ((~II27402));
assign g26143 = ((~g8296))|((~g14725))|((~g25438))|((~g25405));
assign g30294 = ((~g13483)&(~g29990));
assign g13415 = ((~II20544));
assign II13104 = ((~g2));
assign g24255 = ((~II31445));
assign II33321 = ((~g24442));
assign g12853 = ((~g8894));
assign g25453 = (g6142&g24763);
assign g24610 = (g23533&g23521);
assign g5628 = ((~g300));
assign g28795 = ((~g28485)&(~g28015));
assign II31808 = ((~g23675));
assign g7139 = ((~g1481));
assign g27925 = ((~g16276)&(~g27661));
assign g4501 = ((~g822));
assign g29573 = (g28803&g29398);
assign g24607 = ((~II32193));
assign g27964 = ((~g16400)&(~g27680));
assign g17654 = (g4486&g15332);
assign g18820 = ((~g13738)&(~g11922));
assign II30203 = ((~g22717));
assign g10330 = (g5556&g2504);
assign g12890 = ((~g8468)&(~g8489)&(~g8505));
assign II37304 = ((~g27802))|((~II37303));
assign g10009 = (g3254&g4211);
assign g15046 = (g4142&g13161);
assign II34800 = ((~g26229));
assign II40303 = ((~g30487));
assign g22425 = ((~II28969));
assign II36069 = ((~g27493));
assign g21246 = ((~g19984)&(~g5929));
assign II35092 = ((~g26669));
assign g10455 = (g3650&g1953);
assign g16861 = ((~g15829)&(~g13032));
assign II39393 = ((~g15971))|((~II39391));
assign g29469 = (g29345&g19511);
assign II16286 = ((~g7265));
assign g9660 = (g3410&g3948);
assign g13077 = ((~g9822))|((~g7230));
assign g7861 = ((~g1316));
assign g14048 = ((~g11915));
assign II37950 = ((~g28556));
assign II28218 = ((~g14194))|((~II28217));
assign II23258 = ((~g14205))|((~II23256));
assign g3618 = ((~II13207));
assign g18940 = ((~g15647));
assign g4584 = ((~g2779));
assign g11262 = ((~II18191))|((~II18192));
assign g11878 = ((~g11114));
assign g30255 = ((~g16263)&(~g30089));
assign g17795 = (g4725&g15443);
assign g28789 = ((~g28477)&(~g27985));
assign g19063 = (g18679&g14910&g13687&g16254);
assign II40423 = ((~g30579));
assign g13516 = (g6045&g12295);
assign g28441 = (g28133&g9257);
assign II37635 = ((~g28390));
assign g19075 = ((~II25258));
assign g20637 = ((~II27228));
assign II30779 = ((~g22080));
assign g30534 = ((~II40182));
assign g4964 = ((~g2090));
assign g12191 = ((~g8382));
assign g28076 = ((~II36673));
assign g5956 = ((~g204));
assign g17208 = ((~g13576));
assign g5199 = ((~II13801));
assign II22990 = ((~g14321))|((~II22988));
assign g29763 = ((~g16438)&(~g29626));
assign g6623 = ((~g1890));
assign II23133 = ((~g13901))|((~II23131));
assign g18829 = ((~g15222));
assign II36417 = ((~g27462));
assign II15599 = ((~g3566));
assign g26699 = ((~II34704));
assign g11687 = ((~g9117)&(~g9122)&(~g9126));
assign II29083 = ((~g21790));
assign g27202 = ((~II35443));
assign II13140 = ((~g36));
assign II14920 = ((~g1312));
assign II23766 = ((~g13550));
assign g13900 = (g7619&g12821);
assign g12651 = ((~II19771));
assign g6776 = ((~g1230));
assign II14831 = ((~g1517));
assign g16063 = ((~g12804));
assign g22079 = ((~g21343)&(~g19623));
assign g19599 = (g3928&g17348);
assign g8296 = ((~g3649));
assign g7522 = ((~g2917));
assign g10605 = (g3462&g5235);
assign g19168 = ((~II25371));
assign g29512 = ((~II38866));
assign II36289 = ((~g27565))|((~g15923));
assign g19662 = (g646&g18824);
assign g6056 = ((~II14547));
assign g23484 = (g18221&g22681);
assign g18852 = ((~g13815)&(~g12012));
assign g28018 = ((~II36527));
assign g30080 = (g29829&g10996);
assign gbuf218 = (g3040);
assign g29109 = ((~g28654)&(~g17001));
assign g11126 = ((~II18040));
assign II26627 = (g18744&g18772&g18796);
assign g27209 = ((~II35464));
assign g12794 = ((~II19855));
assign g27145 = ((~II35334));
assign g10907 = ((~II17780));
assign II31195 = ((~g22578));
assign g10363 = (g6643&g4746);
assign g9387 = ((~II16590));
assign II18521 = ((~g9449));
assign g9669 = ((~g5552));
assign g24485 = ((~g23625)&(~g22556));
assign g25175 = ((~II33003));
assign g23176 = ((~II29981));
assign g4757 = ((~g718));
assign II21404 = ((~g13037));
assign II27225 = ((~g19358));
assign g29462 = ((~II38767));
assign g4418 = ((~g2105));
assign g25475 = (g14148&g25087);
assign II25634 = ((~g65))|((~II25633));
assign g18956 = ((~g15711));
assign g19976 = (g5330&g18371);
assign g30913 = ((~II40991));
assign g9342 = ((~g5972));
assign g13514 = ((~g12711))|((~g3722));
assign g19837 = (g6901&g17799);
assign g20317 = ((~g17321));
assign g10962 = ((~g5979));
assign II35759 = ((~g27121));
assign g13125 = ((~g9676))|((~g6980));
assign g24899 = (g2046&g23867);
assign II23361 = ((~g15759));
assign II18755 = ((~g9629));
assign g23118 = (g20850&g15890);
assign g23516 = ((~II30560));
assign II28671 = ((~g21845));
assign g10597 = (g7488&g5221);
assign g11518 = ((~II18530));
assign II24272 = ((~g6180))|((~II24271));
assign g22454 = ((~g17012)&(~g21891));
assign II28550 = ((~g21432));
assign g24579 = ((~II32133));
assign II20613 = ((~g12437));
assign II16264 = ((~g6713));
assign II33371 = ((~g25015));
assign g26129 = ((~g8287))|((~g14691))|((~g25431))|((~g25395));
assign g4617 = ((~g717));
assign II17759 = ((~g7263));
assign II25752 = ((~g18390))|((~II25750));
assign g23852 = (g19179&g22696);
assign II27267 = ((~g19358));
assign g29460 = ((~II38761));
assign II30578 = ((~g23124));
assign g4797 = ((~g1414));
assign g4724 = ((~g2504));
assign g26318 = (g4737&g25573);
assign g19287 = ((~g16608));
assign g26829 = (g5623&g26209);
assign g28100 = ((~II36732))|((~II36733));
assign g12798 = ((~II19859));
assign g20722 = ((~II27311));
assign g25502 = ((~II33330));
assign II14002 = ((~g276));
assign g15182 = ((~II21479));
assign g23393 = ((~g22526)&(~g21418));
assign g5824 = ((~g1486));
assign g15130 = ((~II21443));
assign g17720 = ((~g15853));
assign g20404 = ((~g17582));
assign g10588 = (g3678&g5196);
assign g15841 = ((~g13331))|((~g12392));
assign g13848 = ((~g11744));
assign g19499 = (g16943&g14922&g14863);
assign g28941 = ((~g28663)&(~g13343));
assign g23254 = ((~II30215));
assign II40465 = ((~g30671));
assign g11594 = ((~II18758));
assign g22836 = ((~II29629));
assign g11524 = ((~II18548));
assign II35824 = ((~g26805));
assign g15825 = ((~g12657))|((~g6783));
assign II33457 = ((~g24451));
assign g8313 = ((~g3897));
assign g11513 = ((~II18515));
assign g5744 = ((~g2195));
assign II32726 = ((~g14514))|((~II32724));
assign II39029 = ((~g29512));
assign II25643 = ((~g749))|((~g18190));
assign g13585 = ((~g11669));
assign II39848 = ((~g30274));
assign g23711 = ((~II30875));
assign g22578 = ((~g21892)&(~g18982));
assign g19081 = ((~II25264));
assign g27561 = (g24038&g27167);
assign g6023 = ((~g1654));
assign II38145 = ((~g29081));
assign II40647 = ((~g30567));
assign g13192 = ((~g9498));
assign g24482 = ((~g24183));
assign g17023 = (g7420&g15440);
assign g19764 = (g4453&g17637);
assign II30531 = ((~g23076));
assign g15694 = ((~g9488))|((~g9277))|((~g12898));
assign g19584 = (g640&g18756);
assign g9264 = ((~g5938));
assign g11881 = ((~g9870)&(~g9953)&(~g10076));
assign II25147 = ((~g18989));
assign g8722 = (g6751&g7830);
assign g13599 = ((~g12886))|((~g3366));
assign II31109 = ((~g22178));
assign II30905 = ((~g22122));
assign g20364 = ((~g17439));
assign II27026 = ((~g19156));
assign II39359 = ((~g29766))|((~g15880));
assign g25055 = ((~g23955))|((~g6945));
assign II33600 = ((~g24463));
assign g28395 = ((~II37334));
assign g27546 = ((~g26769)&(~g24441));
assign g26355 = ((~II34316));
assign gbuf78 = (g1139);
assign g18566 = ((~g14985));
assign II35146 = ((~g26671));
assign g18449 = ((~II24475))|((~II24476));
assign g30463 = ((~II40027));
assign g3993 = ((~II13275));
assign g27628 = ((~g27038))|((~g3618));
assign II32625 = ((~g17927))|((~II32624));
assign g29983 = (g29885&g8344);
assign g6635 = ((~g2364));
assign II32098 = ((~g24181));
assign g12081 = ((~g10287)&(~g10366)&(~g10433));
assign g30121 = ((~II39628));
assign g20414 = ((~g17621));
assign g28691 = ((~II37620));
assign g16106 = (g12308&g10949);
assign II30332 = ((~g22836));
assign II30911 = ((~g22124));
assign g23159 = ((~II29930));
assign g22271 = ((~g20704));
assign g14194 = ((~g11988));
assign II37008 = ((~g28096));
assign g28948 = (g14222&g28648);
assign g22618 = (g21907&g12756);
assign g17540 = (g4175&g16026);
assign g10104 = (g6448&g4340);
assign g30020 = ((~g29539)&(~g29953));
assign g28269 = ((~II37056));
assign g30864 = ((~II40844));
assign g23221 = ((~II30116));
assign g10173 = (g7265&g2486);
assign II26926 = ((~g17303));
assign g17775 = (g4699&g15432);
assign II22163 = ((~g12433));
assign II24306 = ((~g13983))|((~g15274));
assign g24822 = (g12945&g24164);
assign g3957 = ((~g856));
assign II24476 = ((~g14580))|((~II24474));
assign g15093 = (g7869&g12601);
assign g18543 = ((~g15819));
assign g25060 = ((~g23803))|((~g5556));
assign II31793 = ((~g23472));
assign g25669 = ((~II33495));
assign g29612 = ((~g13933)&(~g29256));
assign g29483 = (g21508&g29286);
assign g13031 = (g7879&g10542);
assign II21881 = ((~g13119));
assign II21761 = ((~g13118));
assign g12871 = ((~II19932));
assign g10375 = (g3462&g1131);
assign II13421 = ((~g2867));
assign g22149 = ((~g21419)&(~g19745));
assign g23340 = ((~g23013))|((~g22189));
assign g18844 = ((~g15284));
assign g19167 = ((~g17556)&(~g15320));
assign g15605 = (g5163&g13256);
assign g16311 = (g5869&g11949);
assign g11945 = ((~g11228));
assign g20841 = ((~g14767)&(~g19552));
assign II13478 = ((~g2854));
assign II15445 = ((~g3236));
assign g30350 = ((~II39873));
assign g15145 = ((~II21458));
assign g21385 = ((~g20492)&(~g13289));
assign g13855 = (g7541&g12691);
assign II27218 = ((~g19168));
assign g24524 = ((~g15494)&(~g23865));
assign g5950 = ((~g2583));
assign II28103 = (g17914&g18358&g17993);
assign g9726 = (g6574&g3978);
assign II17649 = ((~g6293));
assign g27701 = ((~II36114));
assign g24283 = ((~II31523));
assign g20897 = ((~g19635)&(~g17463));
assign g10369 = (g6678&g4760);
assign g13676 = (g5434&g12533);
assign g30940 = ((~II41044));
assign II26317 = (g18295&g18205&g18108);
assign g16141 = (g5706&g11826);
assign g18602 = ((~g16213));
assign II37122 = ((~g28069));
assign g4760 = ((~g720));
assign II24186 = ((~g6177))|((~g13958));
assign g12299 = ((~II19469));
assign g19830 = ((~g18886));
assign g18637 = ((~II24752))|((~II24753));
assign II23932 = ((~g16233));
assign g29913 = ((~II39332))|((~II39333));
assign g10887 = ((~II17750));
assign g26344 = (g4824&g25612);
assign g16425 = (g5968&g12102);
assign g10480 = (g7466&g7342&II17429);
assign g23163 = ((~II29942));
assign g24570 = ((~II32116));
assign g20337 = ((~g16712)&(~g16943));
assign II30380 = ((~g22776));
assign II22775 = ((~g14737));
assign II34132 = ((~g25228));
assign g30519 = ((~II40137));
assign g30500 = ((~g14182)&(~g30222));
assign g19252 = (g18725&g9527);
assign II37143 = ((~g28092));
assign II26123 = ((~g17503));
assign g27506 = ((~g26861));
assign g30063 = ((~g29812)&(~g11637));
assign g21844 = (g20222)|(g18645)|(II28365);
assign g14106 = ((~g11947));
assign g27909 = (g13895&g27397);
assign II20132 = (g2892&g2903&g7595&g2908);
assign g20150 = ((~g16560)&(~g16954));
assign g18509 = ((~g14541));
assign g13818 = (g7531&g12597);
assign g11246 = ((~II18172));
assign II30311 = ((~g22747));
assign II30353 = ((~g22873));
assign II24596 = ((~g14139))|((~II24594));
assign g12547 = ((~g8696));
assign II28506 = ((~g21377));
assign g9888 = (g3254&g4098);
assign g8303 = ((~g3677));
assign g21188 = (g20140&g12379);
assign II36060 = ((~g27353));
assign II26999 = ((~g19543));
assign II29641 = ((~g20825));
assign II39825 = ((~g30268));
assign g27579 = ((~g26775)&(~g25192));
assign g20684 = ((~II27275));
assign g21825 = ((~II28360));
assign g8898 = ((~II16172));
assign II28781 = ((~g21331));
assign g5768 = (g1018&g1068);
assign g12783 = ((~II19844));
assign g24247 = (g22551&g11297);
assign g28172 = ((~g27475));
assign II39806 = ((~g30310));
assign II25573 = ((~g18286))|((~II25571));
assign g5684 = ((~g900));
assign II39832 = ((~g30270));
assign g27000 = (g23340&g26568);
assign II16835 = ((~g3494));
assign g25069 = ((~g24014))|((~g7303));
assign g15725 = (g5296&g13293);
assign II35768 = ((~g26941));
assign g14041 = ((~g8873))|((~g12510))|((~g12495));
assign g15797 = ((~g13305)&(~g7143));
assign g5067 = ((~g1420));
assign g20466 = ((~g17865));
assign g24503 = ((~g23747)&(~g22650));
assign g13434 = ((~II20601));
assign g14514 = ((~g12180));
assign II32616 = ((~g18247))|((~II32615));
assign g4310 = ((~g2254));
assign g24420 = ((~II31934));
assign g15962 = ((~g11675));
assign g20250 = ((~g18764));
assign II38440 = ((~g28738));
assign g26748 = ((~II34851));
assign II40188 = ((~g30347));
assign g18934 = ((~g15628));
assign g28461 = ((~g27729)&(~g26787));
assign g19942 = (g14438&g18536&II26396);
assign g5785 = ((~g1683));
assign g12444 = ((~II19608));
assign g13132 = ((~g9968))|((~g7488));
assign g8030 = ((~II15326));
assign g16905 = ((~II22866));
assign g27583 = ((~g26887))|((~g1430));
assign II28557 = ((~g21407));
assign II28966 = ((~g20633));
assign g27022 = (g21996&g26590);
assign g6215 = ((~g978));
assign g10296 = (g6713&g4644);
assign g23156 = ((~II29921));
assign II30329 = ((~g22800));
assign g25242 = ((~g24802)&(~g23630));
assign g29227 = ((~g28986)&(~g28486));
assign II32499 = ((~g18155))|((~II32498));
assign g12273 = (g8172&g8829);
assign II38698 = ((~g29331));
assign II40817 = ((~g30738));
assign II35904 = ((~g27051))|((~g14831));
assign g22547 = ((~g21087));
assign g11202 = ((~II18124));
assign g29655 = ((~II39083));
assign II31835 = ((~g23911));
assign g21577 = ((~II28111));
assign g13274 = ((~g8906)&(~g8939)&(~g8972));
assign II35506 = ((~g26909));
assign g30742 = ((~II40510));
assign g24241 = (g22259&g11228);
assign g27395 = ((~g26989))|((~g5438));
assign g22581 = (g21895&g12699);
assign II22503 = ((~g13598));
assign g5293 = ((~g738));
assign II34421 = ((~g25203));
assign g30722 = ((~II40456));
assign g21685 = ((~g20164))|((~g6232));
assign g22806 = ((~g21615));
assign g13644 = ((~g13215));
assign g26859 = ((~II35021))|((~II35022));
assign II18593 = ((~g9390));
assign g5806 = ((~g249));
assign II24166 = ((~g14768));
assign g9107 = (g5512&g7718);
assign II24053 = ((~g6777))|((~g14286));
assign II14384 = ((~g3218));
assign g25557 = ((~II33385));
assign II13971 = ((~g1757));
assign g30394 = (g30237&g8990);
assign g22038 = ((~g21305)&(~g19565));
assign II37312 = ((~g27897))|((~II37311));
assign g23003 = ((~g21667))|((~g1358));
assign g16656 = ((~II22699));
assign g23950 = ((~g22992)&(~g6707));
assign g8798 = ((~II16002));
assign II33954 = ((~g25343));
assign g28116 = (g27613&g10316);
assign g23894 = (g22971&g9936);
assign g13458 = ((~II20673));
assign g29183 = (g29064&g20739);
assign II13601 = ((~g121));
assign II27949 = ((~g19957));
assign g18688 = (g14811&g14910&g16254&g13756);
assign g26661 = ((~g25337)&(~g17122));
assign g23572 = (g3934&g22448);
assign g26250 = ((~II34204));
assign g20994 = ((~g19808)&(~g17836));
assign II38184 = ((~g28837));
assign g21207 = (g19456&g19430&II27772);
assign g20087 = (g16749&g7574);
assign II21476 = ((~g11672));
assign g11709 = ((~g9676))|((~g3522));
assign g29471 = (g21461&g29266);
assign g13040 = ((~g9822))|((~g7358));
assign II23374 = ((~g15807));
assign g28158 = ((~g27416));
assign II24408 = ((~g6298))|((~II24407));
assign g10262 = (g7265&g4575);
assign II25054 = ((~g14837));
assign g16830 = ((~II22797));
assign II27388 = ((~g19401));
assign g5704 = ((~g219));
assign g27911 = ((~g16170)&(~g27657));
assign g22917 = ((~g21703));
assign g10468 = (g7265&g4997);
assign g7632 = ((~g1000));
assign g16057 = ((~g12794));
assign g25162 = ((~II32964));
assign g21428 = (g9427&g20420);
assign II29177 = ((~g20900));
assign g21721 = ((~g20198))|((~g6369));
assign g20991 = ((~g19804)&(~g17814));
assign g11182 = ((~II18100));
assign g23021 = ((~g21530));
assign g17649 = ((~II23733));
assign II30881 = ((~g22114));
assign g9114 = (g7015&g7739);
assign g27446 = (g18142&g27141);
assign g19825 = ((~II26266));
assign g8778 = (g3650&g8079);
assign g22382 = ((~g14584))|((~g21189))|((~g10735));
assign g25225 = ((~g24773)&(~g23583));
assign g13493 = (g5887&g11613);
assign II36114 = ((~g27522));
assign g24583 = ((~II32143));
assign g25895 = ((~g24939));
assign g27165 = ((~g23484)&(~g26074));
assign g8524 = (g3566&g1636);
assign g21508 = ((~g19987));
assign g21182 = (g20080&g20103);
assign g8820 = ((~II16034));
assign II33999 = ((~g25490));
assign g8529 = (g6838&g2333);
assign II23395 = ((~g15785));
assign II34866 = ((~g26618));
assign g25985 = ((~II33807));
assign g27655 = ((~g26842)&(~g26061));
assign g7425 = ((~II14990));
assign g19615 = (g1378&g18788);
assign II34059 = ((~g25207));
assign g24567 = ((~II32109));
assign g25931 = ((~g24989))|((~g7015));
assign g26325 = (g4746&g25582);
assign g22643 = (g14016&g21505);
assign g29701 = ((~II39157));
assign II26006 = ((~g16866));
assign g17719 = (g2993&g16065);
assign II18378 = ((~g6314));
assign g27970 = (g14238&g27475);
assign II18423 = ((~g5778));
assign g21695 = (g3554&g20517);
assign g4453 = ((~g132));
assign g13249 = ((~g10018));
assign II13745 = ((~g1506));
assign II21644 = ((~g13096));
assign g10413 = (g7488&g4873);
assign g11783 = ((~g10966));
assign g17246 = ((~g16046)&(~g16066));
assign II21435 = ((~g11662));
assign II32181 = ((~g24238));
assign g28288 = ((~II37113));
assign II22318 = ((~g13370))|((~II22316));
assign gbuf191 = (g2455);
assign gbuf166 = (g1900);
assign g17193 = (g7766&g14420);
assign II15645 = ((~g6783));
assign II30239 = ((~g22834));
assign II26407 = ((~g17132));
assign g12600 = ((~g8766));
assign II16159 = ((~g5403));
assign g27062 = (g22093&g26628);
assign g21872 = ((~g19749));
assign g23497 = ((~g22876)&(~g5606));
assign g13837 = (g7556&g12642);
assign g15839 = ((~g12711))|((~g7085));
assign II38272 = ((~g29013));
assign g12981 = ((~g10354)&(~g6890));
assign II36687 = ((~g27318));
assign II31811 = ((~g24055));
assign g19697 = (g653&g18838);
assign g10145 = (g7162&g4383);
assign g14423 = ((~g12120));
assign g10038 = ((~g7772))|((~g3366));
assign g30499 = (g30191&g11435);
assign g15391 = (g4752&g13205);
assign g29261 = (g28867&g8941);
assign II38653 = ((~g29307));
assign g23080 = ((~g21158)&(~g19324)&(~g19347));
assign g16535 = (g15161&g13774&g13805&g13825);
assign g20578 = ((~II27059));
assign g4489 = ((~g730));
assign g27029 = (g23368&g26600);
assign g13703 = (g8018&g11848);
assign g5618 = ((~g3093));
assign g27971 = ((~II36438));
assign g28056 = ((~II36621));
assign II28335 = (g20254)|(g20241)|(g20217);
assign g21263 = ((~g20064)&(~g5992));
assign g15625 = ((~II21878));
assign g20427 = ((~g17670));
assign II20376 = ((~g8569));
assign II28432 = ((~g19335));
assign g19272 = ((~II25567));
assign g9288 = ((~g5363));
assign g4326 = ((~g181));
assign g29409 = ((~g28840)&(~g28389));
assign II24466 = ((~g9453))|((~II24464));
assign g12820 = ((~g8396)&(~g8438)&(~g8466));
assign g12435 = ((~II19587));
assign g29222 = ((~g28958)&(~g28479));
assign g12204 = ((~II19380));
assign II22136 = (g13082&g2912&g7522);
assign g22975 = ((~g21756));
assign g16820 = ((~g15161));
assign II21583 = ((~g13080));
assign g27672 = ((~g26799)&(~g10024));
assign g10473 = (g7303&g5005);
assign g10394 = (g7053&g4829);
assign g18059 = (g5126&g15644);
assign g12022 = ((~g11348));
assign g14092 = ((~g12890));
assign g24122 = ((~g22458));
assign g26559 = ((~g13824)&(~g25287));
assign II31077 = ((~g22882));
assign II32411 = ((~g24037))|((~II32409));
assign g29190 = ((~II38275));
assign g24611 = (g2151&g23940);
assign g5200 = ((~II13804));
assign II32559 = ((~g17927))|((~g24081));
assign g18084 = ((~g14068));
assign g24784 = ((~II32320));
assign g21085 = (g19484&g14158&g19001);
assign g16686 = ((~g14811));
assign g21352 = (g9391&g20350);
assign g30675 = ((~g16416)&(~g30495));
assign g23097 = ((~g17079)&(~g21161));
assign g15650 = (g5132&g12901);
assign II25018 = ((~g14366));
assign g23324 = ((~g22144)&(~g10024));
assign g21141 = (g20178&g12315);
assign g13407 = ((~II20520));
assign II25690 = ((~g753))|((~g17741));
assign g25255 = ((~g24838)&(~g23714));
assign g29127 = ((~g28376)&(~g27779));
assign g30852 = ((~II40808));
assign g6513 = ((~g660));
assign II28515 = ((~g21557));
assign II33157 = ((~g25027));
assign II30679 = ((~g22049));
assign II40498 = ((~g30681));
assign g19733 = (g672&g18855);
assign g16451 = (g5818&g13386);
assign II24459 = ((~g13599));
assign g29371 = ((~g28932));
assign II26996 = ((~g19169));
assign g16444 = (g5981&g12135);
assign g17063 = ((~g14719));
assign g19414 = ((~II25839))|((~II25840));
assign g17979 = ((~II24016))|((~II24017));
assign g9871 = (g7085&g4082);
assign g11644 = ((~g9076)&(~g9092)&(~g9102));
assign g12938 = (g8179&g10096);
assign g12107 = ((~g10312)&(~g10389)&(~g10451));
assign II32709 = ((~g23892))|((~II32708));
assign g5909 = ((~g1630));
assign g13612 = ((~II20836));
assign g26081 = ((~g25470)&(~g25482));
assign g16220 = (g1896&g11879);
assign g8860 = ((~II16110));
assign g23223 = ((~II30122));
assign II19160 = ((~g10549));
assign g24889 = ((~II32616))|((~II32617));
assign g23172 = ((~II29969));
assign g21346 = ((~g20480)&(~g13247));
assign g5641 = ((~g3185));
assign II36963 = ((~g28030));
assign g10481 = ((~g7826));
assign II37602 = ((~g28579));
assign g10469 = (g5556&g5000);
assign II38817 = ((~g29354));
assign g13475 = ((~II20709));
assign g15415 = ((~II21677));
assign g20669 = ((~II27260));
assign g20022 = ((~g17204))|((~g1466));
assign II38136 = ((~g28833));
assign g13609 = (g6141&g12456);
assign g4567 = ((~g2239));
assign g9670 = ((~II16763));
assign II24247 = ((~g16337));
assign g13396 = ((~II20497));
assign g30233 = ((~g30031));
assign g15750 = ((~II21998));
assign II25617 = ((~g1426))|((~II25616));
assign g27356 = (g65&g26987);
assign g19430 = ((~II25866))|((~II25867));
assign g28820 = ((~II37781));
assign II16972 = ((~g3900));
assign g13054 = ((~g9968))|((~g7488));
assign g22683 = ((~II29333));
assign II31817 = ((~g24077));
assign g5837 = ((~g2374));
assign g29438 = ((~II38695));
assign g19182 = ((~II25399));
assign g12267 = ((~g8460));
assign g26925 = ((~g25648))|((~g26327));
assign II25377 = ((~g18743));
assign g26741 = ((~II34830));
assign II30470 = ((~g23117));
assign g23103 = ((~g21682));
assign g8605 = ((~g6887));
assign g20160 = (g18170&g9424);
assign g22707 = (g14177&g21566);
assign II32057 = ((~g23406));
assign g27989 = ((~II36468));
assign g10987 = ((~g6015));
assign g27277 = ((~g27005)&(~g26318));
assign g9073 = (g7195&g1947);
assign g19040 = ((~II25183));
assign g23141 = ((~g21825));
assign g22090 = ((~g21352)&(~g19637));
assign II36330 = ((~g27447));
assign g11530 = ((~II18566));
assign II24634 = ((~g14467))|((~II24632));
assign g9212 = ((~II16486));
assign II18405 = ((~g5720));
assign g16241 = (g5805&g11892);
assign II28190 = ((~g14079))|((~II28189));
assign g5078 = ((~g1955));
assign g23665 = (g17825&g22995);
assign g11425 = ((~II18389));
assign g25708 = ((~g24728)&(~g24509));
assign II27689 = ((~g19070));
assign g22922 = ((~II29712));
assign g23040 = ((~g14378)&(~g14290)&(~g21142));
assign g29632 = ((~II39014));
assign g18717 = (g14863&g14991&g16313&g13797);
assign II16234 = ((~g5420));
assign g29778 = ((~g29479)&(~g29229));
assign II31112 = ((~g22179));
assign g12174 = ((~g8366));
assign g18370 = ((~II24388))|((~II24389));
assign g25938 = ((~g25129)&(~g17065));
assign II24125 = ((~g14201))|((~II24123));
assign g24296 = ((~II31562));
assign g27084 = (g23388&g26641);
assign g10206 = (g3410&g4498);
assign g24321 = ((~II31637));
assign g20934 = ((~g19714)&(~g17617));
assign g20564 = ((~II27017));
assign II23466 = ((~g15838));
assign g25153 = ((~II32937));
assign g4295 = ((~g2226));
assign g11769 = ((~II18943));
assign g26589 = ((~g25606));
assign II39148 = ((~g29616));
assign g4204 = ((~g3188));
assign g19208 = ((~II25445));
assign g26163 = (g1365&g25939);
assign g22666 = (g21825&g20014);
assign II26777 = ((~g17222));
assign g24265 = ((~II31469));
assign g17527 = (g4254&g15198);
assign gbuf94 = (g1069);
assign g30759 = (g30588&g22360);
assign g13914 = (g7626&g12851);
assign II33573 = ((~g24513));
assign g4737 = ((~g376));
assign g20343 = ((~g16856)&(~g13703));
assign II21677 = ((~g13075));
assign g21758 = (g7607&g20045);
assign g11918 = ((~g11176));
assign II33624 = ((~g24466));
assign g27741 = ((~g27407)&(~g26966));
assign g21688 = ((~g20198))|((~g6519));
assign g21762 = ((~g19471)&(~g18004)&(~g14194));
assign gbuf133 = (g1669);
assign g30972 = ((~II41090));
assign g15311 = ((~II21580));
assign g25553 = (g14385&g25105);
assign g22656 = ((~II29274));
assign g20115 = (g16804&g3139);
assign g17685 = ((~II23769));
assign g26470 = (g5252&g25830);
assign g27248 = (g27037&g16733);
assign g24799 = (g12916&g24149);
assign g21328 = (g9187&g20327);
assign g9647 = (g6678&g3942);
assign g10533 = (g7303&g5118);
assign g28499 = ((~g26027)&(~g27725));
assign g8397 = ((~II15599));
assign g26001 = ((~II33855));
assign g22162 = ((~g21438)&(~g19770));
assign g21879 = ((~g18419))|((~g19250))|((~g19263));
assign g29199 = ((~g28892)&(~g28448));
assign g16002 = ((~g12604));
assign g16596 = ((~II22651));
assign II23553 = ((~g13525));
assign g17445 = ((~g16250));
assign g25773 = ((~II33608));
assign g15802 = (g8253&g13352);
assign g15761 = ((~g12611))|((~g6519));
assign g20585 = ((~II27080));
assign II34099 = ((~g25219));
assign II34806 = ((~g26230));
assign II40044 = ((~g30256));
assign II15967 = ((~g3494));
assign II16776 = ((~g3618));
assign g17517 = ((~II23605));
assign g25490 = (g24759)|(g23146);
assign g28474 = (g18226&g27965);
assign g10380 = (g6751&g1282);
assign II34821 = ((~g26314));
assign g24092 = ((~g22020)&(~g20840));
assign g5071 = ((~II13745));
assign g26405 = (g5050&g25717);
assign g10591 = (g3806&g5207);
assign g11002 = ((~II17907));
assign II14668 = ((~g3232));
assign gbuf148 = (g1712);
assign II28447 = ((~g19369));
assign g20106 = (g18261&g3167);
assign II37968 = ((~g28529));
assign II22028 = (g13004&g3018&g7549);
assign g9534 = (g7772&g6135&g538);
assign g5928 = ((~g270));
assign g14079 = ((~g11935));
assign g7751 = ((~g2479));
assign g22235 = (g21726&g12163);
assign g24270 = ((~II31484));
assign II29462 = ((~g21001));
assign II38491 = ((~g28767));
assign g22714 = (g14207&g21573);
assign g29644 = ((~II39050));
assign g7772 = ((~g659));
assign II18725 = ((~g8977));
assign II13501 = ((~g789));
assign g29793 = (g29491&g11063);
assign g17171 = ((~II23218))|((~II23219));
assign gbuf86 = (g1029);
assign g25020 = ((~g23923))|((~g6643));
assign g15951 = ((~g12711))|((~g6838));
assign g24229 = (g22232&g11105);
assign II16881 = ((~g3998))|((~II16879));
assign g26479 = (g5275&g25847);
assign II37062 = ((~g28040));
assign g30661 = ((~g16345)&(~g30467));
assign g29809 = ((~II39279));
assign g20216 = (g16736&g16943&g16712);
assign g5033 = ((~g608));
assign g19324 = (g16895&g16575&g14186);
assign g3999 = ((~g3204));
assign g27175 = ((~g26075)&(~g25342));
assign g16120 = ((~g10952)&(~g6161)&(~g12507));
assign II35994 = ((~g15074))|((~II35992));
assign g10108 = (g6486&g569);
assign g21689 = ((~II28218))|((~II28219));
assign g19417 = ((~g16591));
assign g25995 = ((~II33837));
assign g16566 = ((~II22631))|((~II22632));
assign II14416 = ((~g3222));
assign II36264 = ((~g27621));
assign II36527 = ((~g27524));
assign II38656 = ((~g29315));
assign II16024 = ((~g7591));
assign g23939 = (g18509&g23095);
assign g8612 = (g3338&g6908);
assign g22526 = (g1332&g21867);
assign g23638 = (g4197&g22543);
assign g24923 = ((~II32669))|((~II32670));
assign II41044 = ((~g30928));
assign g12519 = ((~II19689));
assign II39154 = ((~g29582));
assign II14934 = ((~g2003));
assign g22205 = (g16223)|(g20866);
assign II18857 = ((~g10891));
assign II31165 = ((~g22194));
assign g6707 = ((~g666));
assign g15021 = ((~II21381));
assign g13480 = (g6018&g12197);
assign g28457 = (g26131&g28168);
assign g30399 = ((~g30116)&(~g30123));
assign g27861 = ((~II36330));
assign g16321 = (g1898&g11954);
assign g19467 = ((~g16719));
assign II40673 = ((~g30639));
assign g26039 = (g25668&g19523);
assign g11176 = ((~II18094));
assign g28450 = (g17993&g27932);
assign g4656 = ((~g1393));
assign g11291 = ((~II18241));
assign g5708 = ((~g303));
assign g27078 = ((~g4632)&(~g26084));
assign II24214 = ((~g14033))|((~II24213));
assign g12434 = ((~g10929));
assign II21730 = ((~g13089));
assign g18547 = (g13677&g13750&II24619);
assign g14360 = ((~g12968));
assign g7465 = ((~g2));
assign g22098 = ((~g21356)&(~g19650));
assign II18473 = ((~g8839));
assign g21075 = ((~g19930)&(~g18246));
assign g25221 = ((~g24767)&(~g23577));
assign g7875 = ((~II15184))|((~II15185));
assign II28351 = (g19111)|(g19108)|(g19102);
assign g8655 = ((~II15847));
assign II38229 = ((~g28950));
assign g27233 = ((~II35536));
assign g7823 = ((~g2396));
assign II18707 = ((~g8665));
assign II34172 = ((~g25239));
assign II34839 = ((~g26495));
assign g6153 = ((~II14665));
assign g16629 = ((~g15981)&(~g15971)&(~g15952));
assign g10890 = ((~II17759));
assign II24071 = ((~g14747));
assign II32596 = ((~g18014))|((~II32595));
assign g20623 = ((~II27194));
assign II37569 = ((~g28498));
assign g20289 = ((~g17259));
assign g15828 = (g7877&g13398);
assign g8774 = (g6751&g7958);
assign g9747 = (g6838&g3987);
assign g30825 = ((~II40727));
assign g10066 = (g5512&g4283);
assign g7792 = ((~g1703));
assign II36450 = ((~g27485));
assign g26560 = ((~g25281)&(~g24559));
assign g20378 = ((~g17487));
assign II40197 = ((~g30371));
assign g26024 = (g25301&g21102);
assign g29073 = ((~II38032));
assign g15283 = (g4548&g13191);
assign g27159 = ((~g26442));
assign g13623 = (g5428&g12472);
assign II38391 = ((~g28730));
assign II38804 = ((~g29353));
assign II19602 = ((~g8940));
assign II34671 = ((~g26192));
assign II19455 = ((~g10606));
assign g26668 = (g25283&g21076);
assign II38032 = ((~g28344));
assign g21283 = (g20357&g16820&g16781);
assign g27688 = ((~II36075));
assign II35123 = ((~g26107))|((~g26096));
assign g29163 = ((~II38232));
assign gbuf214 = (g2632);
assign g23821 = ((~II31043));
assign g7259 = ((~g2046));
assign II36302 = ((~g27379))|((~II36300));
assign g26549 = ((~g25421));
assign II39331 = ((~g29705))|((~g29751));
assign II18344 = ((~g7015));
assign II25731 = ((~g758))|((~g18091));
assign g16994 = (g7819&g15323);
assign gbuf47 = (g395);
assign g10549 = ((~g7999));
assign g22864 = ((~II29656));
assign II37917 = ((~g28328));
assign II31826 = ((~g23895));
assign g19455 = ((~g17177));
assign g27790 = (g5875&g27376);
assign g27194 = ((~II35419));
assign g24853 = (g12974&g24180);
assign g15615 = ((~II21871));
assign g12181 = ((~II19360));
assign g21323 = (g9471&g20322);
assign g13206 = ((~g9644));
assign g16433 = ((~g13066));
assign II24415 = ((~g14053))|((~g15366));
assign g27387 = ((~II35727));
assign g21360 = (g9507&g20361);
assign g5860 = ((~g924));
assign g29278 = ((~II38405));
assign g24788 = (g15618&g24140);
assign g30895 = ((~II40937));
assign g25458 = ((~II33282));
assign g13223 = ((~g9816));
assign g20398 = ((~g17560));
assign g28837 = ((~II37804));
assign g26485 = ((~II34449));
assign g25077 = ((~g23414)&(~g22196));
assign g12250 = ((~g10513)&(~g10571)&(~g10615));
assign g11148 = ((~II18064));
assign II35953 = ((~g26824));
assign g16262 = (g1204&g11904);
assign g17573 = ((~II23661));
assign II22545 = ((~g15018));
assign g7303 = ((~II14951));
assign g13146 = ((~g9968))|((~g7426));
assign II24565 = ((~g14472))|((~g9595));
assign g11539 = ((~II18593));
assign g9025 = ((~II16347));
assign g17655 = ((~II23739));
assign g22081 = ((~g21345)&(~g19625));
assign g8626 = (g7195&g7479);
assign g13116 = ((~g9676))|((~g6980));
assign g23120 = (g21819)|(g21814);
assign g25103 = ((~II32829));
assign II23673 = ((~g13539));
assign g15670 = (g5241&g13272);
assign g15356 = (g2020&g12762);
assign g13361 = ((~II20448));
assign g22173 = ((~g21456)&(~g19791));
assign g30950 = (g30932&g20819);
assign g6038 = ((~g2279));
assign II33816 = ((~g25647));
assign g29959 = (g29774&g29035);
assign g19770 = (g4498&g17655);
assign g6288 = ((~g287));
assign g13255 = ((~g10049));
assign II36666 = ((~g27551))|((~g14966));
assign II18259 = ((~g5778));
assign g30989 = ((~II41141));
assign II19631 = ((~g10801));
assign II32588 = ((~g23937))|((~II32586));
assign g7014 = ((~II14882));
assign g13487 = (g5874&g11608);
assign g11637 = (g5918&g8427);
assign g22791 = ((~II29559));
assign II15671 = ((~g3566));
assign g30365 = ((~II39906));
assign g21019 = ((~g19851)&(~g17947));
assign g28715 = (g28414&g22332);
assign g10566 = (g3494&g5156);
assign g19101 = (g18708&g14922&g16313&g13797);
assign II36102 = ((~g27533));
assign g4217 = ((~g354));
assign g26175 = ((~II34077));
assign II18107 = ((~g7875))|((~II18106));
assign g14207 = ((~g12930));
assign II21488 = ((~g11673));
assign II24236 = ((~g9613))|((~II24234));
assign g18825 = ((~g15198));
assign g5886 = ((~II14338));
assign II27005 = ((~g19164));
assign II32970 = ((~g24556));
assign g5639 = ((~g2588));
assign g26794 = (g26143&g16647);
assign g29667 = ((~g29524)&(~g29294));
assign g29235 = (g9453&g28807);
assign g27470 = ((~g26790)&(~g25198));
assign g20187 = (g13805&g13825&II26630);
assign II18097 = ((~g6838));
assign g25050 = ((~g23803))|((~g5556));
assign g3940 = ((~g408));
assign g5793 = ((~g2170));
assign g27875 = ((~g27521)&(~g14677));
assign g8236 = ((~g2219));
assign g22046 = (g21117&g21105&g21096&II28594);
assign g29205 = ((~g15143)&(~g28923));
assign g30309 = ((~II39770));
assign g5550 = ((~II14030));
assign g12239 = ((~II19412));
assign II35053 = ((~g26655));
assign g29292 = ((~g28820));
assign g10613 = (g3494&g1297);
assign g3942 = ((~g699));
assign g17927 = ((~II23976));
assign g23873 = ((~II31133));
assign g15290 = ((~II21566));
assign II16006 = ((~g3878));
assign g29658 = ((~g29574));
assign II40829 = ((~g30815));
assign g26971 = (g23325&g26546);
assign g29026 = ((~g9187))|((~g28512));
assign g28490 = ((~g27240)&(~g27721));
assign II30965 = ((~g22140));
assign g11364 = ((~II18320));
assign II27382 = ((~g19390));
assign g20703 = ((~g20164))|((~g3254));
assign II38841 = ((~g29333))|((~g15981));
assign g24355 = ((~II31739));
assign g20441 = ((~II26874));
assign g26096 = ((~g6068)&(~g24183)&(~g25394));
assign g11209 = ((~II18133));
assign g6443 = ((~g2821));
assign g23127 = (g20858&g15923);
assign g25418 = ((~g24482)&(~g22319));
assign II18662 = ((~g8996));
assign g27991 = (g14360&g27498);
assign g23525 = (g5929&g22787);
assign g19263 = (g17887)|(g17979);
assign g4133 = ((~g848));
assign g21901 = ((~g13552)&(~g19355));
assign g23539 = ((~g22942)&(~g5697));
assign g11309 = ((~II18259));
assign II20547 = ((~g13248));
assign g30953 = (g8605&g30952);
assign II40143 = ((~g30329));
assign g15661 = ((~g11737)&(~g7345));
assign g30034 = ((~II39533))|((~II39534));
assign II30728 = ((~g22065));
assign g8147 = ((~g857));
assign g11891 = ((~g11132));
assign g27518 = ((~II35886));
assign II29336 = ((~g20954));
assign g13572 = ((~II20794));
assign g25755 = ((~II33586));
assign II33408 = ((~g25040));
assign g28832 = ((~II37793));
assign II18746 = ((~g8707));
assign g27308 = ((~g27048)&(~g26387));
assign g24436 = (g14669&g15933&g24134);
assign g30554 = ((~II40242));
assign g25044 = ((~g23955))|((~g6751));
assign g28955 = ((~II37924));
assign g8439 = (g6369&g927);
assign II36721 = ((~g27328));
assign g26333 = (g4772&g25593);
assign g14153 = ((~g12913));
assign g30472 = (g30163&g11300);
assign II13968 = ((~g1078));
assign g28479 = (g18286&g27973);
assign g5132 = ((~g2802));
assign g24728 = ((~g23907)&(~g22788));
assign II25882 = ((~g17914))|((~II25880));
assign g23899 = (g22975&g9962);
assign g11984 = ((~g11287));
assign II39014 = ((~g29535));
assign g29802 = ((~II39258));
assign g10121 = (g3462&g1110);
assign g16814 = ((~II22786));
assign II34143 = ((~g25231));
assign g26385 = ((~II34343));
assign g21963 = ((~II28515));
assign II24502 = ((~g14044))|((~II24500));
assign g11475 = ((~II18441));
assign II25153 = ((~g18995));
assign g26269 = (g4512&g25510);
assign g24975 = ((~g23497))|((~g74));
assign g23629 = ((~II30757));
assign g8089 = ((~II15354));
assign II31715 = ((~g23566));
assign II41141 = ((~g30988));
assign g10943 = ((~II17840));
assign g19300 = ((~II25634))|((~II25635));
assign g19817 = (g2040&g18901);
assign g20936 = ((~g19716)&(~g17619));
assign g20962 = ((~g19758)&(~g17714));
assign g29218 = ((~g15282)&(~g28966));
assign g21856 = (g20284)|(g18655)|(II28380);
assign g21128 = (g19534&g14507&g16560);
assign gbuf97 = (g1084);
assign g26059 = ((~g25422))|((~g25379))|((~g25274));
assign g15235 = (g4437&g13184);
assign g24309 = ((~II31601));
assign g19034 = ((~II25165));
assign II27065 = ((~g19270));
assign II40075 = ((~g30262));
assign g24752 = (g9507&g24106);
assign g21311 = (g9471&g20306);
assign g26294 = ((~II34254));
assign g15464 = ((~II21723));
assign g7574 = ((~g3128));
assign II14766 = ((~g545));
assign g26812 = ((~g15321)&(~g26291));
assign II29383 = ((~g20972));
assign II27537 = ((~g19957));
assign g23409 = (g21533&g22408);
assign g22733 = ((~II29439));
assign g23402 = ((~g18622))|((~g22922));
assign g20290 = ((~g17262));
assign g30389 = (g30233&g8928);
assign g26978 = (g21976&g26551);
assign II40712 = ((~g30652));
assign g30093 = (g29853&g11222);
assign g18611 = ((~II24717))|((~II24718));
assign g30221 = (g30044&g8993);
assign g18806 = ((~g15109));
assign g17635 = (g4322&g16043);
assign g21482 = (g15210&g20446);
assign II28374 = (g20307)|(g18689)|(g18667);
assign g30324 = ((~II39815));
assign g23148 = ((~II29897));
assign g8466 = (g3410&g924);
assign II23941 = ((~g13946))|((~g9293));
assign g18108 = ((~g14537));
assign II38471 = ((~g28758));
assign g24344 = ((~II31706));
assign II33640 = ((~g24467));
assign II25168 = ((~g16877));
assign g19589 = (g8224&g17324);
assign g10432 = (g6486&g4894);
assign g17272 = ((~II23358));
assign II30786 = ((~g22454));
assign II40967 = ((~g30778));
assign g9140 = ((~II16444));
assign g19872 = (g1352&g18928);
assign g16020 = ((~g6200)&(~g12457)&(~g10952));
assign g10876 = ((~II17737));
assign II28271 = ((~g14431))|((~g19515));
assign II15183 = ((~g2975))|((~g2978));
assign II14091 = ((~g2258));
assign II38107 = ((~g28368));
assign g26493 = (g5312&g25862);
assign g28676 = ((~II37575));
assign g26867 = ((~II35043))|((~II35044));
assign g29975 = ((~II39463));
assign g18014 = ((~II24049));
assign g18405 = ((~g14609));
assign II29180 = ((~g20779));
assign g23460 = ((~II30496));
assign g26725 = ((~II34782));
assign g20493 = ((~g18401))|((~g2720));
assign g19925 = (g2059&g18962);
assign g16650 = (g15296&g15366);
assign g20306 = ((~g17294));
assign g9131 = (g6713&g7785);
assign II34241 = ((~g25252));
assign II27056 = ((~g19196));
assign g27569 = ((~II35983));
assign II22283 = ((~g2962))|((~II22282));
assign g30490 = (g30183&g11398);
assign g23622 = (g4136&g22520);
assign g15374 = (g4720&g13203);
assign g18707 = ((~g13636)&(~g11788));
assign II40658 = ((~g30572));
assign g27135 = ((~g26178));
assign g18363 = ((~II24373))|((~II24374));
assign g28583 = ((~II37502));
assign g30402 = ((~g29999)&(~g30129));
assign g11563 = ((~II18665));
assign g23316 = ((~II30401));
assign II19642 = ((~g10793));
assign II37641 = ((~g28375));
assign g20830 = ((~II27419));
assign g13308 = ((~g10273));
assign g24769 = (g9649&g24123);
assign g18789 = ((~g15065));
assign II31748 = ((~g23711));
assign g8812 = ((~II16024));
assign g21092 = (g20124&g14431&g14514);
assign II29715 = ((~g21094));
assign g13028 = ((~g9534))|((~g6678));
assign II16694 = ((~g3462));
assign g5613 = ((~II14069));
assign g21050 = ((~g20513));
assign g8649 = ((~II15839));
assign g22787 = ((~g21199));
assign g20925 = ((~g19708)&(~g17598));
assign g28712 = (g28406&g22276);
assign II39785 = ((~g30124));
assign II39585 = ((~g29941));
assign g10974 = ((~II17875));
assign g26967 = (g6212&g26202);
assign g28554 = ((~g27806));
assign g25176 = ((~II33006));
assign g26994 = (g23331&g26562);
assign g3246 = ((~II13134));
assign g15260 = ((~g12198));
assign II17743 = ((~g8107));
assign g12705 = ((~II19797));
assign g27681 = (g26788&g11456);
assign II36393 = ((~g27572));
assign g30506 = ((~II40098));
assign II31541 = ((~g23500));
assign II16196 = ((~g6116));
assign g24500 = ((~g23740)&(~g22643));
assign g28629 = ((~g27889));
assign II29906 = ((~g21967));
assign g8979 = (g7391&g2568);
assign g7619 = ((~g999));
assign g30412 = ((~II39982));
assign II37002 = ((~g28056));
assign g30466 = ((~II40032));
assign g27344 = ((~g27100)&(~g26478));
assign g19321 = ((~II25691))|((~II25692));
assign g23126 = ((~g17144)&(~g21203));
assign g11788 = (g1240&g8632);
assign g10735 = ((~g4671));
assign g18296 = ((~II24299))|((~II24300));
assign g16848 = ((~II22820));
assign g11532 = ((~II18572));
assign g21345 = (g15096&g20346);
assign g30819 = ((~II40709));
assign g30107 = (g29873&g11382);
assign g4272 = ((~g1542));
assign g12040 = ((~g11367));
assign g23464 = ((~II30504));
assign g18900 = ((~g15496));
assign g29179 = ((~g28849)&(~g28405));
assign II31943 = ((~g24000));
assign II26365 = ((~g18626));
assign g30380 = ((~II39945));
assign II14709 = ((~g3229));
assign II30931 = ((~g22129));
assign II33472 = ((~g24499));
assign g30343 = ((~II39856));
assign g19576 = (g8197&g17310);
assign g10439 = (g3462&g4913);
assign g29315 = ((~II38474));
assign g29925 = ((~II39368))|((~II39369));
assign g25609 = ((~II33434));
assign g26229 = ((~II34165));
assign II15190 = ((~g2956))|((~g2959));
assign g4041 = ((~g864));
assign g22066 = ((~g21334)&(~g19604));
assign g20299 = ((~g16665)&(~g16884));
assign g30958 = ((~g30922)&(~g30948));
assign g12941 = ((~g8504)&(~g8519)&(~g8534));
assign g10399 = (g7358&g4842);
assign g16614 = ((~g15962)&(~g15942)&(~g14677));
assign II38662 = ((~g29253));
assign g22843 = ((~g21889));
assign g11957 = ((~g10081)&(~g10172)&(~g10259));
assign g21715 = ((~g20164))|((~g6314));
assign g26673 = (g12431&g25318);
assign II26645 = (g14849&g18728&g13687);
assign II35945 = ((~g27078))|((~II35944));
assign g8878 = ((~II16144));
assign g27690 = ((~II36081));
assign g29537 = ((~II38909));
assign II36969 = ((~g28031));
assign II29536 = ((~g21027));
assign g28759 = ((~g28442)&(~g27935));
assign g4827 = ((~g1816));
assign II19797 = ((~g10147));
assign g15831 = ((~g13313))|((~g12392));
assign II28991 = ((~g20648));
assign II36659 = ((~g27312));
assign g21748 = ((~g20228))|((~g6783));
assign g8868 = (g6751&g1177);
assign g1248 = ((~II13092));
assign g16006 = ((~g12984))|((~g7426));
assign g29038 = ((~g9216))|((~g28567));
assign II27285 = ((~g19420));
assign II15535 = ((~g6519));
assign g25351 = (g24683&g18120);
assign g23119 = (g5904&g21069);
assign II19030 = ((~g8726));
assign g22725 = ((~II29421));
assign g16492 = ((~II22578));
assign g21413 = (g15188&g20405);
assign II38379 = ((~g28845))|((~II38378));
assign g28469 = (g18179&g27952);
assign g24949 = ((~II32704));
assign g16825 = ((~g15855));
assign g8505 = (g3410&g942);
assign II27779 = ((~g20022));
assign g26569 = ((~g13837)&(~g25290));
assign g29141 = ((~II38166));
assign II31445 = ((~g22687));
assign g24641 = ((~g1880))|((~g23394));
assign II37956 = ((~g28584));
assign g21948 = ((~II28470));
assign g25287 = (g24687&g8757);
assign g30510 = ((~II40110));
assign g6485 = ((~II14766));
assign g16384 = (g296&g12024);
assign g20631 = ((~II27218));
assign g17937 = ((~g13983));
assign g17761 = ((~II23836));
assign II17981 = ((~g7976));
assign II13504 = ((~g793));
assign g28024 = ((~II36539));
assign g11527 = ((~II18557));
assign II16357 = ((~g3774));
assign g12647 = ((~II19767));
assign II30504 = ((~g22936));
assign II34860 = ((~g26548));
assign g29196 = (g15022&g28741);
assign g7573 = ((~g3120));
assign g27380 = ((~II35708));
assign g18782 = ((~g13676)&(~g13705));
assign g30761 = (g30621&g20822);
assign II19618 = ((~g10814));
assign g10478 = (g7488&g5018);
assign g13974 = ((~g11872));
assign II23636 = ((~g15851));
assign II18302 = ((~g3254));
assign g22181 = ((~g21486)&(~g19815));
assign g12155 = ((~g10386)&(~g10450)&(~g10514));
assign g7532 = ((~g1471));
assign II15454 = ((~g3239));
assign II25253 = ((~g17124));
assign g16967 = (g7827&g15175);
assign g9661 = (g6519&g3951);
assign g22188 = ((~II28727))|((~II28728));
assign g22223 = (g21921&g12109);
assign g12880 = ((~g8465)&(~g8486)&(~g8502));
assign g23714 = (g4401&g22592);
assign g28216 = ((~II36897));
assign g15032 = ((~g12027));
assign g23543 = ((~II30589));
assign g20566 = ((~II27023));
assign g8908 = ((~II16190));
assign g26234 = (g4343&g25479);
assign g9481 = ((~II16650));
assign II21615 = ((~g13090));
assign g10745 = (g3678&g5382);
assign g4465 = ((~g346));
assign g17429 = ((~g16239)&(~g16288));
assign g22596 = (g20928&g17613);
assign g5960 = ((~g882));
assign g5664 = ((~g65));
assign g20826 = (g5770&g19118);
assign g26652 = ((~g25841));
assign II39919 = ((~g30294));
assign g11973 = ((~g11278));
assign g5388 = ((~II13892));
assign II33385 = ((~g25035));
assign II20640 = ((~g11670));
assign g26018 = ((~II33906));
assign g24400 = ((~II31874));
assign g11138 = ((~II18052));
assign II16438 = ((~g3522));
assign g27431 = ((~g27066))|((~g7265));
assign g21053 = ((~g19901)&(~g18107));
assign g25027 = ((~g24227)&(~g17001));
assign g30390 = (g30229&g8952);
assign II16107 = ((~g5398));
assign II13892 = ((~g3040));
assign g28853 = (g27892&g28624);
assign g8274 = ((~II15490));
assign g26365 = (g4913&g25652);
assign g11934 = ((~g10011)&(~g10104)&(~g10193));
assign g13548 = ((~g12611))|((~g3410));
assign g19919 = ((~II26369));
assign g9734 = ((~II16785));
assign g14238 = ((~g12939));
assign II34971 = ((~g26557));
assign g10670 = (g3806&g5312);
assign g18074 = ((~g14062));
assign g23532 = ((~II30578));
assign g17209 = ((~g8160)&(~g14493));
assign II35485 = ((~g27180));
assign g12538 = ((~g8305))|((~g7265));
assign g23683 = ((~II30841));
assign II27300 = ((~g19390));
assign II40709 = ((~g30651));
assign II26085 = ((~g18085));
assign II38396 = ((~g28727));
assign g13189 = ((~g9468));
assign g17202 = ((~g14737))|((~g14753));
assign g23145 = ((~g21825));
assign g21597 = (g13927&g14268&g19843&II28126);
assign g8388 = ((~II15590));
assign g25121 = ((~II32851));
assign gbuf101 = (g1237);
assign g13530 = ((~g13251));
assign II31152 = ((~g22191));
assign g23448 = ((~II30476));
assign g30768 = ((~II40559))|((~II40560));
assign II33649 = ((~g25063));
assign g8839 = ((~II16071));
assign g25237 = ((~g24793)&(~g23610));
assign g16395 = ((~g13049));
assign g21435 = ((~g20503)&(~g16385));
assign g19621 = (g3987&g17378);
assign II15546 = ((~g6783));
assign g29561 = ((~II38947));
assign g9057 = (g7053&g1945);
assign g25618 = (g7259&g25110);
assign g29934 = ((~II39404));
assign g11958 = ((~g11246));
assign II37074 = ((~g28084));
assign II37280 = ((~g28179));
assign II40691 = ((~g30645));
assign g10452 = (g7015&g4948);
assign II38722 = ((~g29319));
assign g29986 = (g29877&g8366);
assign II16335 = ((~g3618));
assign g11949 = ((~g11234));
assign g8714 = ((~II15918));
assign II36493 = ((~g27266));
assign g16847 = ((~g15095)&(~g12650));
assign g27097 = (g22134&g26650);
assign g11435 = ((~II18399));
assign g26567 = ((~g25543));
assign g4015 = ((~g411));
assign g29456 = ((~II38749));
assign g24293 = ((~II31553));
assign g15220 = ((~g12163));
assign g21340 = (g9737&g20340);
assign g25826 = ((~g24638)&(~g24533));
assign g21953 = ((~II28485));
assign g30871 = ((~II40865));
assign g18325 = ((~g14736))|((~g10082));
assign g28082 = ((~II36687));
assign g10063 = (g6783&g4278);
assign g11404 = ((~II18362));
assign g17167 = (g8009&g15764);
assign g20422 = ((~g17655));
assign g23728 = ((~II30908));
assign g12075 = ((~g11411));
assign g21173 = (g20095&g16575&g16523);
assign g5064 = ((~g1409));
assign II28123 = ((~g19987));
assign II33662 = ((~g24532));
assign g26340 = (g4783&g25602);
assign g4905 = ((~g723));
assign g28166 = ((~g27451));
assign g29280 = ((~g28791));
assign g13529 = ((~g12611))|((~g3410));
assign II38851 = ((~g29169));
assign II23029 = ((~g14221))|((~II23027));
assign g15755 = (g8178&g13309);
assign II18375 = ((~g3254));
assign g5859 = ((~g805));
assign g10520 = (g3650&g1973);
assign gbuf99 = (g1018);
assign g28244 = ((~II36981));
assign g8573 = (g7085&g2282);
assign g19354 = ((~g14768))|((~g8605))|((~g17157));
assign g21316 = ((~g20460)&(~g16111));
assign g26941 = ((~g25835))|((~g26417))|((~g25798));
assign II24263 = ((~g14342))|((~g9232));
assign II38857 = ((~g29172));
assign g23922 = ((~g4456)&(~g22985));
assign g17716 = (g4584&g15382);
assign g22607 = (g13946&g21458);
assign II13101 = ((~g1));
assign g21887 = ((~g13519)&(~g19289));
assign g27089 = (g22118&g26646);
assign g24263 = ((~II31463));
assign g11999 = ((~g10166)&(~g10250)&(~g10319));
assign g26025 = ((~g25392)&(~g17193));
assign g27312 = ((~g27054)&(~g26397));
assign g23604 = (g4064&g22494);
assign g4101 = ((~g161));
assign g23309 = ((~II30380));
assign g20940 = ((~g19723)&(~g17633));
assign g4541 = ((~g1735));
assign g26681 = ((~II34650));
assign g21377 = ((~II27920));
assign g19309 = ((~II25660));
assign g22985 = ((~g21618)&(~g21049));
assign II14778 = ((~g823));
assign g6912 = ((~II14860));
assign g21293 = ((~II27838));
assign g26896 = ((~II35095));
assign g19931 = (g14637&g14139&II26383);
assign g17366 = ((~II23454));
assign II24124 = ((~g6290))|((~II24123));
assign g11579 = ((~II18713));
assign g28782 = ((~g15304)&(~g28475));
assign g28334 = (g27842&g20793);
assign g15898 = ((~g12657))|((~g6574));
assign g24779 = (g9569&g24131);
assign II14249 = ((~g3216));
assign II37134 = ((~g28107));
assign II19307 = ((~g8726));
assign g15807 = ((~g12611))|((~g6369));
assign g19812 = (g4674&g17755);
assign g4003 = ((~g158));
assign g18221 = ((~g14747));
assign II30803 = ((~g22089));
assign g16895 = ((~g13589));
assign g29325 = ((~II38496));
assign II25283 = ((~g17086));
assign g26763 = (g14691&g26516);
assign II28464 = ((~g21024));
assign g22004 = (g978&g21202);
assign g13285 = ((~g10189));
assign g22669 = ((~II29301));
assign g26188 = (g2753&g25945);
assign II27116 = ((~g19762));
assign g18618 = ((~II24726))|((~II24727));
assign g28748 = ((~g28435)&(~g27924));
assign g4928 = ((~g1279));
assign g10305 = (g6980&g4662);
assign g30089 = (g29835&g11160);
assign g10227 = (g3618&g4545);
assign g5238 = ((~g1270));
assign g30565 = ((~II40275));
assign g13049 = ((~g10851));
assign g25505 = (g6707&g25094);
assign g7153 = ((~g480));
assign g11627 = ((~g9063)&(~g9077)&(~g9093));
assign g11896 = ((~g9903)&(~g10036)&(~g10112));
assign II36996 = ((~g28055));
assign g11582 = ((~II18722));
assign II36272 = ((~g15890))|((~II36270));
assign g19546 = ((~II25971));
assign g24590 = (g23486&g23478);
assign g8252 = ((~g2861));
assign g24676 = (g13568&g24115);
assign g29404 = ((~II38599));
assign g10867 = ((~g5850));
assign II41050 = ((~g30938));
assign g18667 = (g14863&g14991&g13724&g16313);
assign II24608 = ((~g16006));
assign g20138 = (g18261&g9756);
assign g12454 = ((~II19634));
assign g30315 = ((~II39788));
assign II28741 = ((~g21890))|((~g13530));
assign g18063 = ((~g15660));
assign g23847 = ((~II31091));
assign g26556 = ((~g25510));
assign g11967 = (g7967&g8711);
assign II30236 = ((~g22866));
assign g22144 = ((~g21410)&(~g19730));
assign g5751 = ((~g52));
assign g4632 = ((~g996));
assign g17551 = ((~II23639));
assign II24916 = ((~g14776));
assign II37032 = ((~g28037));
assign g25144 = ((~II32910));
assign g19046 = ((~II25201));
assign g17947 = (g4964&g15563);
assign g25257 = ((~g24841)&(~g23722));
assign g15756 = ((~g13313))|((~g12354));
assign g8761 = (g7195&g8156);
assign g5903 = ((~II14357));
assign II18620 = ((~g11385));
assign g20356 = ((~g17425));
assign II29936 = ((~g22582));
assign g22742 = ((~II29462));
assign II38875 = ((~g29184));
assign gbuf67 = (g558);
assign g10574 = ((~g8013));
assign g3677 = ((~g1880));
assign II15304 = ((~g1855));
assign g8911 = ((~g5114));
assign g20805 = ((~g20255))|((~g3722));
assign g24460 = ((~g23748))|((~g3618));
assign II30594 = ((~g22025));
assign II30401 = ((~g22444));
assign g19161 = (g17207&g8627);
assign g27365 = (g1439&g27036);
assign II31619 = ((~g23597));
assign gbuf196 = (g2400);
assign g29759 = ((~g16379)&(~g29622));
assign g25065 = ((~g23984))|((~g7053));
assign gbuf11 = (g2833);
assign g16133 = (g6444&g11817);
assign g24104 = ((~g22422));
assign g4486 = ((~g714));
assign g9521 = (g3254&g8200);
assign g18753 = (g14936&g15080&g16371&g13825);
assign g27215 = ((~II35482));
assign g9463 = (g6369&g8144);
assign g14464 = ((~g12153));
assign g21817 = (g20219)|(g20187)|(II28346);
assign II37179 = ((~g27784));
assign g18491 = ((~II24531))|((~II24532));
assign g6166 = ((~II14675));
assign g19771 = (g4501&g17658);
assign II33888 = ((~g25817));
assign g7265 = ((~II14945));
assign g27005 = (g23331&g26578);
assign II35079 = ((~g26664));
assign g30966 = ((~g30956));
assign g17912 = (g4908&g15537);
assign g11778 = ((~g10949));
assign II24389 = ((~g13974))|((~II24387));
assign g22342 = ((~g21172))|((~g21249))|((~g21156));
assign g10996 = ((~II17901));
assign II30894 = ((~g22117));
assign g29689 = ((~II39121));
assign g11770 = ((~g10932));
assign g17384 = ((~II23472));
assign g21541 = ((~II28076));
assign g24864 = ((~g23473));
assign g4203 = ((~g20));
assign g12148 = ((~g8333));
assign II29927 = ((~g23105));
assign g29063 = ((~g28326)&(~g28329));
assign g29382 = ((~g28993));
assign g5118 = ((~g2653));
assign g23046 = ((~g21128)&(~g19282));
assign II23115 = ((~g13848))|((~II23113));
assign g20622 = ((~II27191));
assign g12415 = ((~II19563));
assign g22935 = ((~g21903)&(~g7466));
assign g25304 = (g24704&g8798);
assign g26414 = (g5078&g25735);
assign g24425 = ((~II31949));
assign II33517 = ((~g25060));
assign g27017 = (g23340&g26585);
assign g25430 = ((~g24616));
assign g4185 = ((~g2228));
assign g24638 = ((~g23673)&(~g22595));
assign g29994 = (g29889&g8418);
assign g25678 = ((~II33504));
assign g27053 = (g23368&g26619);
assign g26259 = (g4471&g25499);
assign g6783 = ((~II14834));
assign II17670 = ((~g6441));
assign II31832 = ((~g23896));
assign g25204 = ((~g24745)&(~g23547));
assign g29905 = ((~g29688));
assign g22061 = ((~g21326)&(~g19593));
assign g26895 = ((~II35092));
assign II18524 = ((~g9640));
assign g19660 = (g633&g18822);
assign g27397 = ((~II35737));
assign II38701 = ((~g29401));
assign g20985 = ((~II27534));
assign g26979 = (g23331&g26552);
assign g16211 = (g1203&g11871);
assign gbuf31 = (g280);
assign g19914 = (g3018&g18958);
assign II24950 = ((~g14922));
assign g16644 = ((~II22687));
assign g22362 = ((~g14529))|((~g21169))|((~g10714));
assign II37494 = ((~g27766));
assign II23806 = ((~g14062))|((~g9150));
assign g23153 = ((~II29912));
assign II18787 = ((~g10910));
assign II16747 = ((~g6643));
assign g27742 = ((~g27409)&(~g26967));
assign II23457 = ((~g15836));
assign g23181 = ((~II29996));
assign g11281 = ((~II18229));
assign g18107 = (g5167&g15675);
assign g25915 = ((~g24951));
assign g11837 = ((~g11045));
assign g20050 = (g18070&g3161);
assign g28636 = ((~g28191)&(~g17065));
assign g28279 = ((~II37086));
assign II31454 = ((~g23727));
assign g11703 = ((~g9132)&(~g9137)&(~g9139));
assign II31763 = ((~g23745));
assign II33495 = ((~g24455));
assign II36808 = ((~g27354));
assign g21162 = (g20038&g20062);
assign g30850 = ((~II40802));
assign g11598 = ((~II18770));
assign g28487 = (g18390&g27999);
assign g23592 = (g17640&g22986);
assign g11459 = ((~II18423));
assign g23094 = ((~II29841));
assign II17910 = ((~g7532));
assign g27289 = ((~g27023)&(~g26344));
assign g24875 = ((~II32568))|((~II32569));
assign g10261 = (g7265&g2495);
assign II32320 = ((~g23979));
assign g6448 = ((~II14763));
assign g27355 = (g61&g26837);
assign g19564 = (g8123&g17272);
assign g18526 = ((~g14559));
assign II22952 = ((~g15210))|((~g14206));
assign g29548 = (g28784&g29383);
assign g29966 = (g29755&g12004);
assign g7459 = ((~g2356));
assign g9083 = (g5556&g7664);
assign g21422 = (g15210&g20412);
assign g24415 = ((~II31919));
assign g5851 = ((~g74));
assign II35021 = ((~g26110))|((~II35020));
assign g18977 = ((~g15797))|((~g3006));
assign II17816 = ((~g7346));
assign g29329 = (g29096&g29002);
assign II32346 = ((~g17815))|((~II32345));
assign g29840 = ((~g29669));
assign g13878 = (g7610&g12782);
assign II31127 = ((~g22183));
assign g25980 = (g24663&g21928);
assign g4590 = ((~II13538));
assign g29119 = ((~II38125));
assign g5716 = ((~g753));
assign g13873 = ((~g12698));
assign II29613 = ((~g21053));
assign g17116 = (g7649&g14008);
assign g5705 = ((~g225));
assign g11914 = ((~g9939)&(~g10073)&(~g10164));
assign g19500 = (g14991)|(g16739);
assign II18943 = ((~g9149));
assign g20502 = (g17566&g11973);
assign II29360 = ((~g21796));
assign g5651 = ((~g758));
assign gbuf112 = (g1214);
assign g23300 = ((~II30353));
assign g28669 = (g27897&g22233);
assign II39930 = ((~g30297));
assign g13055 = (g7471&g7570&II20100);
assign g27048 = (g22009&g26614);
assign g15019 = ((~II21377));
assign II18204 = ((~g7975))|((~g4202));
assign g9891 = (g3254&g4107);
assign II24743 = ((~g6167))|((~g14486));
assign g30869 = ((~II40859));
assign g29529 = (g29199&g29370);
assign g17507 = ((~g16298)&(~g13318));
assign II18777 = ((~g9050));
assign g30844 = ((~II40784));
assign g29535 = ((~II38905));
assign II16876 = ((~g7303));
assign g19347 = (g16895&g16546&g14273);
assign g10014 = (g5438&g429);
assign II18566 = ((~g8825));
assign g13934 = ((~g8587))|((~g12478));
assign g9922 = (g3566&g4156);
assign g4945 = ((~g1742));
assign g17393 = (g3941&g16005);
assign II33659 = ((~g24469));
assign g12034 = ((~g10200)&(~g10286)&(~g10365));
assign g28894 = ((~II37863));
assign II38408 = ((~g28721));
assign g29607 = (g29193&g11056);
assign g25315 = ((~II33145));
assign g3235 = ((~II13101));
assign g6430 = ((~g1670));
assign g3243 = ((~II13125));
assign g23505 = ((~g22885))|((~g14584))|((~g10735));
assign II13128 = ((~g26));
assign g29410 = ((~II38613));
assign g13464 = ((~II20691));
assign g13632 = ((~II20858));
assign g23315 = ((~II30398));
assign II36123 = ((~g27540));
assign g20738 = ((~g20198))|((~g3410));
assign g9591 = ((~II16700));
assign g11591 = ((~II18749));
assign g19688 = (g2766&g18834);
assign g26531 = ((~g25974)&(~g17065));
assign g7607 = ((~g2924));
assign g20679 = ((~II27270));
assign g12863 = ((~II19924));
assign g20457 = ((~II26892));
assign II19628 = ((~g10784));
assign g24055 = ((~II31274));
assign g24644 = (g17203&g24115);
assign g13600 = ((~II20820));
assign II31655 = ((~g23739));
assign II19105 = ((~g8726));
assign g28962 = (g14292&g28650);
assign g13881 = ((~g11789));
assign II30525 = ((~g23067));
assign g29264 = (g28867&g8997);
assign g11589 = ((~II18743));
assign g26070 = ((~II33968));
assign g16770 = ((~g14991));
assign g30919 = (g30786&g22297);
assign II33434 = ((~g25025));
assign g8406 = (g6783&g1597);
assign II16156 = ((~g5438));
assign g4415 = ((~g2085));
assign II30763 = ((~g22076));
assign g21789 = (g19128)|(g16913)|(g14811);
assign g18874 = ((~g15412));
assign g22231 = ((~g21666)&(~g19971));
assign gbuf189 = (g2442);
assign g10289 = (g6912&g4614);
assign g15744 = ((~II21992));
assign g24507 = ((~g15391)&(~g23824));
assign II17060 = ((~g6637))|((~II17059));
assign g15784 = ((~g12565))|((~g6232));
assign g18952 = ((~II24992));
assign II27095 = ((~g19185));
assign g22182 = ((~g21487)&(~g19821));
assign g30539 = ((~II40197));
assign g20145 = (g14776&g18670&g16142&g16189);
assign g25184 = (g24694&g20735);
assign g12996 = ((~g9038));
assign g25179 = ((~II33013));
assign g30929 = ((~g30728)&(~g30736));
assign II24061 = ((~g14207))|((~g9326));
assign g27717 = ((~II36162));
assign II31290 = ((~g22269));
assign g20012 = (g16804&g3135);
assign II16120 = ((~g5400));
assign g18832 = ((~g15231));
assign g28265 = ((~II37044));
assign g9794 = (g6980&g4052);
assign g26113 = ((~g25426)&(~g22319));
assign g19213 = (g18030)|(g18115);
assign g30071 = ((~g29834)&(~g29839));
assign g9762 = (g3254&g4009);
assign g6641 = ((~g113));
assign II39913 = ((~g30292));
assign g23972 = (g2903&g23115);
assign g7898 = ((~g3057));
assign g22307 = ((~g20772));
assign g23677 = ((~II30829));
assign g25372 = ((~g24997)&(~g5689));
assign g20554 = ((~g18587));
assign g20016 = ((~II26458));
assign g17080 = ((~II23066))|((~II23067));
assign g21996 = ((~g19268))|((~g21159))|((~g19312));
assign II18329 = ((~g5720));
assign g18867 = ((~g13835)&(~g12070));
assign g29726 = ((~g29503));
assign g22628 = ((~II29226));
assign g10556 = (g3338&g611);
assign g21195 = (g20212&g12385);
assign g15845 = ((~g12565))|((~g6314));
assign g30935 = ((~g30760)&(~g30762));
assign g5213 = ((~g2656));
assign g19705 = ((~II26134));
assign g24835 = ((~II32439));
assign g8958 = ((~II16264));
assign g20297 = ((~g17275));
assign II37273 = ((~g28179));
assign g24212 = ((~g16987)&(~g22244));
assign II34114 = ((~g25958));
assign g21397 = (g9342&g20393);
assign g13958 = ((~g11863));
assign g30687 = ((~g13479)&(~g30345));
assign g16170 = (g3616&g11842);
assign g21009 = ((~g19839)&(~g17900));
assign g26196 = ((~II34114));
assign g9905 = (g3410&g4127);
assign II26340 = ((~g17025));
assign g8843 = ((~II16079));
assign II23742 = ((~g15888));
assign g26539 = ((~g25463));
assign g5879 = ((~g2306));
assign g14107 = ((~g12893));
assign g25361 = ((~g24837));
assign g8723 = (g6945&g8071);
assign II29951 = ((~g22584));
assign g13120 = ((~g9822))|((~g7358));
assign g21628 = ((~II28159));
assign II17070 = ((~g7528));
assign g19767 = (g666&g18872);
assign g11712 = ((~g9968))|((~g3834));
assign g12913 = ((~g8487)&(~g8503)&(~g8518));
assign g23024 = ((~g21537));
assign g30455 = ((~g13953)&(~g30216));
assign g18246 = (g5286&g15747);
assign g18805 = ((~g15106));
assign g18985 = ((~II25047));
assign g18586 = ((~II24678))|((~II24679));
assign g8414 = ((~II15616));
assign g27113 = (g1248)|(g1245)|(g26534);
assign g16356 = (g1206&g11989);
assign g11225 = ((~II18151));
assign g29131 = ((~II38136));
assign g22613 = ((~II29197));
assign II37863 = ((~g28529));
assign g5921 = ((~g2582));
assign II18810 = ((~g10813));
assign g5686 = ((~II14134));
assign g20324 = ((~g17333));
assign g30461 = (g30163&g11234);
assign g25954 = ((~g22806))|((~g24517));
assign g23797 = (g23128)|(g21938);
assign g25437 = ((~g24627));
assign g30653 = ((~g16289)&(~g30454));
assign gbuf151 = (g1893);
assign II36621 = ((~g27301));
assign g8763 = ((~II15955));
assign g11826 = ((~g11028));
assign g19780 = (g4532&g17679);
assign II35731 = ((~g26892));
assign g30064 = ((~g29813)&(~g13506));
assign g7337 = ((~g2190));
assign g13791 = ((~g12444));
assign g6204 = ((~g289));
assign g22992 = ((~g21636))|((~g672));
assign g24457 = ((~g23923))|((~g3338));
assign g27096 = (g23388&g26649);
assign g10372 = (g3462&g4769);
assign g16236 = ((~g12935));
assign II28988 = ((~g20874));
assign II37170 = ((~g28126));
assign II23173 = ((~g13881))|((~II23171));
assign g13455 = ((~II20664));
assign g6894 = ((~g2362));
assign II29465 = ((~g21002));
assign g24454 = ((~g23955))|((~g3494));
assign g22125 = ((~g21381)&(~g19695));
assign g26758 = (g16614&g26521&g13637);
assign II21888 = ((~g13120));
assign g25347 = ((~g24817));
assign II16344 = ((~g5556));
assign II29116 = ((~g20882));
assign II15478 = ((~g3247));
assign g16693 = ((~g15981)&(~g14737)&(~g15952));
assign II24077 = ((~g14414))|((~II24076));
assign g14960 = ((~II21361));
assign II20328 = ((~g10817));
assign II27355 = ((~g19335));
assign g28121 = ((~II36792));
assign g23031 = ((~g21550));
assign g30680 = ((~g16443)&(~g30327));
assign II14066 = ((~g1564));
assign g18921 = ((~g15569));
assign II28143 = ((~g19957));
assign g30878 = ((~II40886));
assign g5999 = ((~g2342));
assign g8544 = (g7085&g2336);
assign g19259 = ((~II25528));
assign g19712 = (g4269&g17534);
assign g9752 = ((~II16796));
assign g6177 = ((~g633));
assign g29546 = ((~II38924));
assign g22633 = (g20956&g17710);
assign II23242 = ((~g9737))|((~g13882));
assign g13168 = ((~g9306));
assign g13441 = ((~II20622));
assign II17483 = ((~g3900));
assign II15696 = ((~g3722));
assign g19244 = (g18458)|(g18514);
assign II18043 = ((~g7976));
assign g9146 = ((~II16450));
assign II18295 = ((~g6314));
assign II34668 = ((~g26210));
assign g11853 = ((~g11066));
assign g19693 = (g4208&g17490);
assign g6131 = ((~II14644));
assign II40979 = ((~g30800));
assign g17155 = (g7535&g15737);
assign g10787 = ((~II17632));
assign g26841 = ((~II34986));
assign g30694 = ((~g13505)&(~g30367));
assign II40627 = ((~g30602))|((~g30594));
assign II30660 = ((~g22043));
assign g7527 = ((~g3018));
assign g13582 = ((~g12290));
assign II27032 = ((~g19189));
assign g18237 = ((~g14514));
assign II23020 = ((~g14032))|((~II23018));
assign g16456 = (g1677&g12160);
assign II21321 = ((~g11758));
assign g20913 = ((~g19669)&(~g17530));
assign g23483 = (g22945&g8847);
assign g18826 = ((~g15201));
assign g25294 = (g24687&g8775);
assign II25562 = ((~g17724))|((~II25560));
assign g12209 = ((~g8397));
assign g5870 = ((~g1621));
assign II40694 = ((~g30646));
assign g30546 = ((~II40218));
assign g16640 = ((~II22683));
assign g19011 = ((~II25096));
assign g22737 = ((~II29451));
assign g26140 = ((~g24183)&(~g25430));
assign g24627 = ((~g1186))|((~g23387));
assign g5342 = ((~g2691));
assign II29945 = ((~g22583));
assign II24758 = (g14936&g15080&g16325);
assign II13134 = ((~g30));
assign g25340 = ((~g21235))|((~g14618))|((~g10754))|((~g24610));
assign g12325 = ((~g8494));
assign g30922 = (g30788&g22315);
assign g15454 = ((~g9232))|((~g9150))|((~g12780));
assign g27935 = (g4251&g27437);
assign g13824 = (g7533&g12598);
assign g15540 = ((~g9310))|((~g9174))|((~g12819));
assign g6193 = ((~II14688));
assign g5473 = ((~II14009));
assign g30143 = ((~g30012));
assign g12061 = ((~g10255)&(~g10323)&(~g10401));
assign g6062 = ((~II14565));
assign g25009 = ((~g23644))|((~g6448));
assign g24163 = ((~g22560));
assign g4347 = ((~g438));
assign g18147 = ((~II24157))|((~II24158));
assign g14355 = ((~g12082));
assign g7084 = ((~II14897));
assign g17056 = (g7953&g15525);
assign II23658 = ((~g14885));
assign g27549 = ((~g26765)&(~g19093));
assign g19386 = ((~II25801))|((~II25802));
assign II36521 = ((~g27274));
assign II40584 = ((~g30704));
assign II27215 = ((~g19158));
assign II21374 = ((~g12424));
assign g20891 = ((~g19626)&(~g17447));
assign II19271 = ((~g10500));
assign II23392 = ((~g13476));
assign g22777 = ((~g21796));
assign g22762 = ((~II29506));
assign II31787 = ((~g23531));
assign g24313 = ((~II31613));
assign g8974 = ((~II16286));
assign g26105 = ((~II34002));
assign g30586 = ((~II40310));
assign II21949 = ((~g11725));
assign II38241 = ((~g28832));
assign g22112 = ((~g21370)&(~g19670));
assign g18090 = ((~II24103))|((~II24104));
assign g24209 = ((~g16984)&(~g22238));
assign g15096 = ((~g11800));
assign g5257 = ((~g2099));
assign g27390 = ((~g26989))|((~g6448));
assign g17604 = ((~II23692));
assign II34189 = ((~g25242));
assign g25385 = ((~g24801));
assign g5867 = ((~g1491));
assign g22847 = ((~g21643));
assign g20604 = ((~II27137));
assign g10889 = ((~II17756));
assign g21895 = ((~g19945));
assign II16562 = ((~g6000));
assign g13501 = ((~g12711))|((~g3722));
assign II15879 = ((~g3678));
assign II35428 = ((~g26953));
assign II20622 = ((~g12543));
assign g29447 = ((~II38722));
assign g24284 = ((~II31526));
assign g30118 = (g29889&g11468);
assign g21370 = (g9326&g20369);
assign II20365 = ((~g9084));
assign g24818 = (g12916&g24162);
assign g4692 = ((~g1819));
assign g29454 = ((~II38743));
assign g20373 = ((~g17479));
assign g18835 = ((~g13788)&(~g11966));
assign II27695 = (g19318&g19300&g19286);
assign g29677 = ((~g29543)&(~g29321));
assign g20403 = ((~g17579));
assign g17224 = ((~g16004)&(~g16009));
assign g7622 = ((~g1852));
assign g11940 = ((~g10044)&(~g10119)&(~g10208));
assign g30048 = ((~g29920));
assign g27226 = ((~II35515));
assign g10801 = ((~g5688)&(~g5729)&(~g5767));
assign g9139 = (g3618&g7809);
assign II35863 = ((~g26811));
assign g11519 = ((~II18533));
assign II16138 = ((~g7053));
assign g6908 = ((~g484));
assign g14316 = ((~g12060));
assign II15909 = ((~g5745));
assign g27769 = ((~g27570)&(~g27111));
assign g16301 = (g5862&g11943);
assign g25869 = ((~II33717));
assign g8160 = ((~g2241));
assign g9063 = (g5438&g7629);
assign II24300 = ((~g14028))|((~II24298));
assign II31901 = ((~g23847));
assign II29687 = ((~g21770));
assign II23929 = ((~g15151));
assign g7993 = ((~g145));
assign g30524 = ((~II40152));
assign g7976 = ((~II15288));
assign g15537 = ((~II21796));
assign g22295 = ((~g20749));
assign g22016 = ((~g21576))|((~g21605));
assign g13318 = ((~II20379));
assign g19920 = (g1372&g18961);
assign g29297 = ((~II38434));
assign g23069 = ((~g21619));
assign g9932 = ((~II16936));
assign g24813 = (g21825&g23905);
assign II13575 = ((~g1476));
assign g30734 = ((~II40490));
assign g20039 = (g5372&g18523);
assign g19853 = (g2046&g18921);
assign II17869 = ((~g7534));
assign g16404 = ((~g13079));
assign g24844 = ((~II32469))|((~II32470));
assign II33330 = ((~g25019));
assign g26617 = ((~g25694));
assign II24507 = ((~g15999));
assign g19453 = ((~II25889))|((~II25890));
assign g22753 = ((~g21184));
assign g25945 = ((~g24827));
assign g30971 = ((~g30970));
assign g23138 = (g20866&g15952);
assign II29550 = ((~g21032));
assign g28057 = (g27599&g10049);
assign g10276 = ((~II17238));
assign g17259 = ((~II23345));
assign g28610 = ((~g27843));
assign g21593 = (g16498&g19484&g14071);
assign g19728 = (g4332&g17560);
assign II30383 = ((~g22803));
assign II38650 = ((~g29314));
assign g13245 = ((~g10779))|((~g7901));
assign g28050 = (g27590&g10018);
assign g19791 = (g4567&g17707);
assign II24235 = ((~g14222))|((~II24234));
assign g19009 = ((~II25092));
assign g20955 = ((~g19754)&(~g17697));
assign II40230 = ((~g30362));
assign g19286 = ((~II25596))|((~II25597));
assign g10103 = (g3254&g4335);
assign g10446 = (g3522&g4930);
assign II32487 = ((~g23400));
assign g29606 = ((~g13878)&(~g29248));
assign g25263 = ((~g24874)&(~g17838));
assign g25167 = ((~II32979));
assign g21179 = (g19534)|(g16602)|(g14423);
assign II40113 = ((~g30368));
assign II28482 = ((~g21376));
assign g30884 = ((~II40904));
assign g9341 = ((~II16562));
assign g16486 = ((~II22560));
assign II34395 = ((~g25929));
assign g12744 = ((~II19808));
assign g12232 = ((~g10474)&(~g10534)&(~g10594));
assign g28115 = ((~II36772));
assign g5626 = ((~g121));
assign g24142 = ((~g22500));
assign g16253 = (g5814&g11900);
assign g3462 = ((~II13186));
assign g23152 = ((~II29909));
assign g29161 = ((~II38226));
assign II20556 = ((~g12435));
assign g8499 = (g6838&g2315);
assign g15409 = ((~g12285));
assign g30060 = ((~g29970)&(~g11612));
assign g16884 = ((~g13589));
assign g26217 = ((~g25963)&(~g13320));
assign II40051 = ((~g30257));
assign g5243 = ((~g1408));
assign II35095 = ((~g26670));
assign II35341 = ((~g26120));
assign g20760 = ((~II27349));
assign g23434 = (g22831&g19640);
assign g30134 = ((~g30010));
assign II39035 = ((~g29544));
assign g13425 = ((~II20574));
assign g30711 = ((~II40423));
assign g13451 = ((~II20652));
assign g10797 = ((~g5678)&(~g5710)&(~g5757));
assign g23287 = ((~II30314));
assign g29306 = ((~II38453));
assign g17236 = ((~g16033)&(~g16051));
assign II37400 = ((~g28200));
assign g5385 = ((~g2813));
assign g6897 = ((~g1486));
assign g5438 = ((~II14002));
assign g9323 = ((~II16552));
assign g29399 = ((~g28834)&(~g28378));
assign II16779 = ((~g7015));
assign II30059 = ((~g22620));
assign g19284 = (g18063&g3111);
assign g10094 = (g7426&g4318);
assign g4474 = ((~g435));
assign II24662 = ((~g13621));
assign g23168 = ((~II29957));
assign g23471 = (g18105&g22645);
assign g21415 = ((~II27958));
assign g26551 = ((~g25496));
assign g27529 = ((~g4456)&(~g26873));
assign g26290 = (g4598&g25530);
assign g16367 = (g1899&g11998);
assign g13834 = (g7336&g12599);
assign g13124 = ((~g8613)&(~g8625)&(~g8631));
assign II34776 = ((~g26277));
assign g20407 = ((~g17591));
assign g20581 = ((~II27068));
assign g22825 = ((~II29606));
assign g5507 = ((~g3155));
assign g20652 = ((~II27243));
assign II25899 = ((~g18226))|((~II25897));
assign g11774 = ((~g10937));
assign g15679 = ((~g12385));
assign g11921 = ((~g11185));
assign g19578 = ((~g16884));
assign g23828 = ((~II31056));
assign g28070 = ((~II36653));
assign g8209 = ((~g832));
assign g15177 = ((~g12339));
assign g27231 = ((~II35530));
assign II36507 = ((~g27270));
assign g17228 = ((~g16016)&(~g16029));
assign II18411 = ((~g3566));
assign II39083 = ((~g29519));
assign g8700 = ((~II15902));
assign g23311 = ((~II30386));
assign g27754 = ((~g27446)&(~g26985));
assign II20305 = ((~g9050));
assign II25702 = ((~g18297))|((~II25700));
assign g19550 = ((~II25977));
assign II33260 = ((~g24909));
assign g25247 = ((~g24811)&(~g23638));
assign II19937 = (g9507&g9427&g9356&g9293);
assign II35043 = ((~g26151))|((~II35042));
assign g21791 = ((~g20255))|((~g6838));
assign g20969 = ((~g19768)&(~g15402));
assign g29990 = (g29885&g8397);
assign II35364 = ((~g26304));
assign g6216 = ((~g2066));
assign g24749 = (g15540&g24102);
assign II13950 = ((~g1063));
assign II39020 = ((~g29499));
assign g24554 = (g19977&g18124&g23415);
assign g15545 = (g5056&g13237);
assign II31736 = ((~g23628));
assign g13142 = ((~g9822))|((~g7230));
assign g11063 = ((~II17981));
assign g12362 = ((~g10866));
assign II30476 = ((~g22876));
assign g15426 = ((~II21688));
assign g12858 = ((~g8448)&(~g8473)&(~g8491));
assign g30798 = ((~g16134)&(~g30697));
assign g5114 = ((~g2599));
assign g27892 = ((~g27546)&(~g14711));
assign g19656 = (g4104&g17439);
assign g23943 = ((~II31205));
assign g21573 = ((~II28107));
assign g11552 = ((~II18632));
assign g23415 = ((~g23084));
assign g24476 = ((~g23477)&(~g20127));
assign II21691 = ((~g13078));
assign g5816 = (g1024&g1070);
assign g23786 = ((~II31000));
assign g29372 = ((~g28937));
assign g9102 = (g3306&g7703);
assign g24079 = ((~II31302));
assign g27050 = (g23381&g26617);
assign g28226 = ((~II36927));
assign g22729 = ((~II29429));
assign g19224 = (g18514)|(g18561);
assign g15161 = ((~g12327));
assign g13546 = ((~g12711))|((~g3722));
assign g8971 = ((~II16279));
assign g25218 = ((~g24760)&(~g23571));
assign g22274 = ((~g20708));
assign II23009 = ((~g9203))|((~II23008));
assign g4424 = ((~g2234));
assign g29946 = (g29778&g28906);
assign g23735 = (g22949&g9450);
assign g30195 = ((~g30025));
assign II40317 = ((~g30338));
assign g28751 = ((~II37712));
assign II32677 = ((~g23823))|((~g14165));
assign g4441 = ((~g2774));
assign g9497 = (g6838&g8161);
assign II17798 = ((~g8031));
assign g25514 = (g24488&g20443);
assign II18280 = ((~g7970))|((~g7923));
assign g4868 = ((~g2507));
assign g16013 = ((~g12692));
assign II33396 = ((~g24447));
assign gbuf209 = (g2556);
assign g27573 = ((~g26773)&(~g25188));
assign g11798 = ((~g10867));
assign II34794 = ((~g26125));
assign II41138 = ((~g30971));
assign g5899 = ((~g809));
assign g15765 = (g5333&g13324);
assign g20665 = (g4985&g19081);
assign g7953 = ((~g487));
assign II28027 = ((~g20067));
assign g29979 = ((~II39475));
assign g28331 = (g27802&g22307);
assign g24515 = ((~g23802)&(~g22686));
assign II16507 = ((~g6448));
assign II29591 = ((~g21047));
assign II38214 = ((~g29101));
assign gbuf62 = (g481);
assign g19779 = (g4529&g17676);
assign g22484 = ((~II29030));
assign g10459 = (g7053&g1976);
assign g5362 = ((~g2817));
assign g11421 = (g6232&g222);
assign II29700 = ((~g20700));
assign g15942 = ((~g11666));
assign g24499 = ((~g15325)&(~g23778));
assign g22837 = ((~II29632));
assign g16111 = (g5551&g13215);
assign II22444 = ((~g1900));
assign g20485 = ((~II26934));
assign g20902 = ((~g19661)&(~g17509));
assign g26850 = ((~II35003));
assign g15821 = ((~g12565))|((~g6314));
assign II28789 = ((~g21878));
assign g20081 = (g5385&g18587);
assign g8492 = (g6783&g1624);
assign g15043 = ((~II21398));
assign II16611 = ((~g6000));
assign g18670 = ((~g14797));
assign g22722 = (g2734&g21586);
assign g10542 = ((~II17483));
assign g28148 = ((~g27658)&(~g17100));
assign g17378 = ((~II23466));
assign g23376 = ((~g18435))|((~g22812));
assign g22566 = (g2026&g21872);
assign II14993 = ((~g2697));
assign II18281 = ((~g7970))|((~II18280));
assign g24381 = ((~II31817));
assign II15610 = ((~g3566));
assign g25723 = ((~II33551));
assign g28296 = ((~II37137));
assign g29559 = (g26045&g29390);
assign g20783 = ((~II27372));
assign g21809 = (g19135)|(g19641)|(g16712);
assign II30648 = ((~g22040));
assign g23565 = (g6146&g22437);
assign g20501 = ((~g18334));
assign g24001 = ((~II31235));
assign g25797 = ((~II33636));
assign g25272 = ((~g24905)&(~g18061));
assign II29445 = ((~g20995));
assign g23748 = ((~II30948));
assign g4444 = ((~g2776));
assign g18814 = ((~g15148));
assign II25664 = ((~g2120))|((~g18474));
assign g25155 = ((~II32943));
assign g21225 = ((~g19132));
assign g10640 = (g3806&g2676);
assign g28307 = ((~II37170));
assign g3900 = ((~II13246));
assign g12522 = ((~g8662));
assign g21867 = ((~g19705));
assign g28043 = ((~II36582));
assign II36761 = ((~g27338));
assign g21027 = ((~g19862)&(~g17967));
assign II25001 = ((~g14244));
assign g3997 = ((~g45));
assign g28096 = ((~II36721));
assign g18910 = ((~g15531));
assign g29698 = ((~II39148));
assign II23225 = ((~g9649))|((~g14090));
assign g22055 = ((~g21320)&(~g19587));
assign g8568 = ((~g6230));
assign g21337 = (g9471&g20334);
assign g18654 = (g15065&g16266&g16360);
assign g21899 = (g19323&g11749);
assign II32461 = ((~g18247))|((~II32460));
assign g21307 = (g9453&g20302);
assign g25403 = ((~g24854));
assign II34068 = ((~g25211));
assign II19753 = ((~g9229));
assign II19374 = ((~g10500));
assign g17020 = ((~II22989))|((~II22990));
assign g27543 = ((~II35933));
assign g30291 = ((~g16460)&(~g29987));
assign g30298 = ((~g13496)&(~g29995));
assign g9067 = ((~g5789));
assign g16559 = ((~II22626));
assign II22789 = ((~g14711));
assign g4269 = ((~g1540));
assign g17288 = ((~II23374));
assign g12431 = ((~g8580)&(~g10730));
assign II32898 = ((~g24856));
assign II32835 = ((~g24072));
assign II35799 = ((~g27130));
assign g15493 = ((~g12321));
assign g11804 = ((~g10995));
assign g22996 = ((~g21449));
assign g15766 = ((~II22014));
assign II16931 = (g5830&g6024&g5070&g5071);
assign g23419 = (g22755&g19577);
assign II38898 = ((~g29194));
assign g28799 = ((~II37760));
assign g30777 = ((~II40597));
assign g16448 = (g5984&g12148);
assign g19144 = ((~g17268)&(~g14884));
assign g14233 = ((~g10773))|((~g12527));
assign g29659 = ((~g29571));
assign g24928 = ((~II32678))|((~II32679));
assign g17217 = ((~g13605));
assign g29950 = (g29788&g28937);
assign II30365 = ((~g22664));
assign g30980 = ((~II41114));
assign g22768 = ((~II29522));
assign g22799 = ((~II29579));
assign g26704 = ((~II34719));
assign g5597 = ((~g1200));
assign g29821 = (g29731&g20746);
assign II32267 = ((~g23936))|((~II32265));
assign g17799 = ((~II23874));
assign II35524 = ((~g27166));
assign g30745 = ((~II40515));
assign g17807 = ((~II23879))|((~II23880));
assign II26690 = (g18744&g18772&g16325);
assign II40206 = ((~g30450));
assign II18287 = ((~g8256))|((~g8102));
assign g19164 = ((~II25365));
assign g21911 = (g19350&g11749);
assign g27811 = ((~g6087)&(~g27632)&(~g25404));
assign g27968 = (g4575&g27472);
assign g15440 = ((~g12302));
assign II24361 = ((~g6157))|((~g14525));
assign II16552 = ((~g6713));
assign g13395 = (g5844&g11475);
assign g23016 = ((~g21518));
assign g12002 = ((~g11318));
assign II21494 = ((~g13061));
assign II31694 = ((~g24064));
assign g24535 = ((~g15562)&(~g23894));
assign II34274 = ((~g25256));
assign g25421 = ((~II33249));
assign II40736 = ((~g30660));
assign g28045 = ((~II36588));
assign g27316 = ((~g27058)&(~g26406));
assign g24251 = ((~g22903));
assign g13091 = ((~g9676))|((~g7162));
assign II36981 = ((~g28074));
assign g11652 = ((~II18838));
assign g21242 = ((~g19455)&(~g17168));
assign g18379 = ((~g14390));
assign g5590 = ((~g3158));
assign II24694 = ((~g6146))|((~g14374));
assign II23198 = ((~g9569))|((~g14176));
assign g9005 = ((~II16325));
assign g8178 = ((~g3052));
assign II30302 = ((~g22724));
assign g5056 = ((~g1288));
assign II23605 = ((~g15847));
assign g16335 = (g2591&g11963);
assign g15424 = (g4828&g13211);
assign g10199 = (g6486&g4476);
assign g13411 = ((~II20532));
assign II27164 = ((~g20418));
assign g29105 = ((~II38104));
assign g5827 = (g1712&g1762);
assign II25831 = ((~g18314))|((~II25829));
assign g7990 = ((~g143));
assign g20728 = ((~g20255))|((~g3722));
assign II32424 = ((~g24046))|((~II32422));
assign g23290 = ((~II30323));
assign g25637 = ((~II33460));
assign II22902 = ((~g14000))|((~II22900));
assign g29247 = ((~II38348));
assign g10497 = (g6912&g5038);
assign II15517 = ((~g8089));
assign g23495 = ((~g10694))|((~g14442))|((~g22316));
assign II23066 = ((~g9277))|((~II23065));
assign g26767 = (g26087&g22287);
assign II16624 = ((~g3306));
assign g19855 = (g18131&g16129);
assign g26751 = ((~II34860));
assign g22286 = ((~g20732));
assign g8706 = (g7195&g7888);
assign g27290 = ((~g27024)&(~g26348));
assign g23671 = (g4275&g22560);
assign g15868 = ((~g12611))|((~g6519));
assign II23842 = ((~g15055));
assign g29173 = ((~g28847)&(~g28402));
assign g17029 = ((~g14685));
assign II27369 = ((~g19457));
assign g17462 = (g4147&g15133);
assign g10705 = ((~g3554))|((~g6980));
assign g26304 = ((~g25978)&(~g16451));
assign g16970 = (g7354&g15221);
assign g3494 = ((~II13190));
assign g8424 = ((~II15626));
assign g28916 = ((~II37885));
assign g8432 = (g6314&g243);
assign g13647 = ((~II20873));
assign g23774 = ((~II30976));
assign g24064 = ((~II31282));
assign g15991 = ((~g12548));
assign g17555 = (g4318&g15240);
assign g17131 = ((~II23143))|((~II23144));
assign g26695 = ((~II34692));
assign g7703 = ((~g320));
assign g11035 = ((~II17948));
assign II36758 = ((~g27337));
assign II36557 = ((~g27284));
assign g21183 = ((~g20192)&(~g20221));
assign II39062 = ((~g29504));
assign g7582 = ((~g2185));
assign II22730 = ((~g14691));
assign II29159 = ((~g20896));
assign II31631 = ((~g23662));
assign g13552 = ((~g13299));
assign II21955 = ((~g13144));
assign g26938 = ((~g25725))|((~g26374));
assign II33128 = ((~g24975));
assign g12935 = ((~II19986));
assign g16843 = ((~II22813));
assign g30644 = ((~g16218)&(~g30442));
assign II23233 = ((~g9711))|((~g14291));
assign g4142 = ((~g1098));
assign II31913 = ((~g23468));
assign II14957 = ((~g2827));
assign g23783 = ((~II30991));
assign g28346 = ((~g15546)&(~g28035));
assign II26276 = ((~g16861));
assign g21738 = ((~g19444)&(~g17893)&(~g14079));
assign g28379 = (g27868&g19390&g19369);
assign g21773 = (g3866&g19078);
assign II39788 = ((~g30125));
assign g17613 = ((~II23701));
assign II30335 = ((~g22801));
assign II33593 = ((~g24445));
assign g20609 = ((~II27152));
assign g26641 = ((~g25790));
assign II20571 = ((~g13341));
assign g10035 = (g3366&g4225);
assign g23478 = ((~g22809))|((~g14442))|((~g10694));
assign g29240 = (g9613&g28820);
assign g11902 = ((~g9911)&(~g10047)&(~g10121));
assign II30245 = ((~g22899));
assign g4885 = ((~g448));
assign II23575 = ((~g15843));
assign g21752 = ((~g19110));
assign g5187 = ((~g2096));
assign g28448 = (g17974&g27928);
assign g23878 = (g22975&g9880);
assign II30953 = ((~g22916))|((~II30952));
assign g27735 = ((~g27394)&(~g26961));
assign g17135 = (g7638&g15698);
assign g21868 = ((~g18302))|((~g19214))|((~g19224));
assign g29812 = (g29762&g12223);
assign g29095 = ((~II38080));
assign g29273 = ((~II38396));
assign II18148 = ((~g6369));
assign g7964 = ((~g2938));
assign g10511 = (g3522&g5058);
assign g18256 = (g5289&g15750);
assign g22515 = (g13873&g21382);
assign II29070 = ((~g20707));
assign II24514 = ((~g9342))|((~II24512));
assign g21062 = ((~g19912)&(~g18154));
assign g9588 = ((~II16697));
assign g8347 = ((~II15549));
assign g25148 = ((~II32922));
assign g20600 = ((~II27125));
assign g30961 = ((~g30925)&(~g30951));
assign g25270 = ((~g24898)&(~g18023));
assign g28842 = ((~II37814))|((~II37815));
assign g29909 = (g29735&g19420&g19401);
assign II16479 = ((~g5438));
assign II32646 = ((~g18155))|((~II32645));
assign g19607 = ((~g16910));
assign g22198 = ((~g19924)&(~g21650));
assign II25135 = ((~g16506));
assign g27186 = ((~II35399));
assign II22631 = ((~g13507))|((~II22630));
assign g20837 = ((~II27426));
assign g29330 = (g29038&g29010);
assign g18919 = ((~g15563));
assign g30702 = ((~g14006)&(~g30390));
assign g30847 = ((~II40793));
assign g18926 = ((~g15596));
assign g11504 = ((~II18488));
assign II33700 = ((~g24474));
assign g15622 = ((~g12370));
assign gbuf57 = (g572);
assign g19056 = ((~II25231));
assign II29429 = ((~g20990));
assign g26733 = ((~II34806));
assign g17175 = ((~II23234))|((~II23235));
assign II26593 = (g14811&g18758&g13687);
assign g10323 = (g7085&g4705);
assign II38767 = ((~g29244));
assign II39779 = ((~g30053));
assign g13944 = (g7141&g12874);
assign gbuf1 = (g2930);
assign g24259 = ((~II31451));
assign g8269 = ((~II15475));
assign II30948 = ((~g22536));
assign g8547 = ((~g3398))|((~g3366));
assign g26043 = ((~g25506)&(~g24870));
assign g20280 = (g13677&g16243&II26695);
assign g6017 = ((~g888));
assign g4313 = ((~g2483));
assign g21861 = ((~g19657));
assign g23454 = ((~II30486));
assign II15369 = ((~g3129));
assign g4963 = ((~g1976));
assign II23661 = ((~g16085));
assign g10403 = (g3722&g4857);
assign g13991 = ((~g11881));
assign II15168 = ((~g2981))|((~II15167));
assign g16292 = (g294&g11932);
assign g26054 = (g25944&g21099);
assign II39323 = ((~g29721))|((~g29713));
assign g22115 = ((~g21373)&(~g19677));
assign g9010 = ((~II16332));
assign II24553 = ((~g6163))|((~g14537));
assign g15971 = ((~g11678));
assign g18995 = ((~II25071));
assign g9368 = ((~II16578));
assign g30497 = ((~II40083));
assign g4705 = ((~g2207));
assign g15375 = (g4724&g13204);
assign g8135 = ((~g172));
assign g20380 = ((~g17493));
assign g19905 = (g2066&g18950);
assign II24007 = ((~g15814))|((~II24005));
assign g29031 = ((~g28319)&(~g28324));
assign g28248 = ((~II36993));
assign II18271 = ((~g6838));
assign g30332 = ((~II39835));
assign g3937 = ((~g178));
assign g13336 = ((~II20407));
assign g22264 = (g21766&g12253);
assign g17752 = (g4656&g15412);
assign g24735 = ((~II32251));
assign II31511 = ((~g23640));
assign g8528 = (g7085&g2327);
assign g29930 = ((~II39385))|((~II39386));
assign II15015 = ((~g2700));
assign g28639 = ((~g27919));
assign g16102 = (g6905&g11795);
assign g23836 = ((~II31068));
assign g27331 = ((~g27083)&(~g26445));
assign g13539 = ((~g12611))|((~g3410));
assign g22879 = ((~g21870))|((~g21866))|((~g21862));
assign II24016 = ((~g13907))|((~II24015));
assign g26779 = ((~g26367))|((~g3462));
assign II30922 = ((~g22126));
assign g22268 = ((~g20697));
assign g30814 = ((~II40694));
assign g24012 = ((~g22887))|((~g14614));
assign g14135 = ((~g11964));
assign II28975 = ((~g21688));
assign g13136 = ((~g9822))|((~g7230));
assign g20944 = ((~g19731)&(~g17652));
assign g13351 = ((~g10416));
assign g4775 = ((~g1085));
assign g12564 = ((~II19736));
assign g27416 = ((~II35756));
assign g19230 = (g16985)|(g16965)|(II25477);
assign II14381 = ((~g3223));
assign g5770 = ((~g992));
assign II35067 = ((~g26659));
assign g13437 = ((~II20610));
assign II31036 = ((~g22941))|((~II31035));
assign g26410 = (g25885)|(g25887);
assign g29146 = ((~II38181));
assign g19626 = (g640&g18805);
assign g24563 = (g18630&g23120&g23415);
assign g7134 = ((~g2727));
assign g26772 = ((~g26320))|((~g3306));
assign g16443 = (g5980&g12134);
assign g9723 = (g6783&g3969);
assign g26808 = ((~g15246)&(~g26262));
assign g29782 = ((~g29482)&(~g29234));
assign g10766 = ((~g6676));
assign g16791 = ((~g15065));
assign g28482 = ((~g27731)&(~g26797));
assign g28241 = ((~II36972));
assign II17907 = ((~g5824));
assign g5414 = ((~II13956));
assign II36577 = ((~g27290));
assign g12128 = (g7916&g8785);
assign II18536 = ((~g11101));
assign g18646 = ((~g16341));
assign g20590 = ((~II27095));
assign g25891 = ((~II33737));
assign II34128 = ((~g25227));
assign g16478 = ((~II22536));
assign g24394 = ((~II31856));
assign g16462 = (g2370&g12177);
assign II29243 = ((~g20921));
assign II18494 = ((~g8821));
assign g18813 = ((~g15145));
assign g17675 = (g4523&g15346);
assign g5919 = (g2412&g2458);
assign g24825 = (g9941&g24166);
assign g18261 = ((~g15719));
assign g10492 = (g3338&g5027);
assign g28410 = ((~g27748)&(~g22344));
assign g11768 = ((~g9367)&(~g9441)&(~g9521));
assign g11922 = (g6431&g8690);
assign g21144 = ((~II27705));
assign g30057 = ((~g29967)&(~g13368));
assign II14083 = ((~g325));
assign g25593 = ((~II33418));
assign g26714 = ((~II34749));
assign g13034 = ((~g9534))|((~g6678));
assign g21782 = ((~g19951));
assign II40928 = ((~g30756));
assign g17713 = (g6890&g16063);
assign g30281 = ((~g16426)&(~g30115));
assign II16549 = ((~g3462));
assign II25192 = ((~g18918));
assign II38160 = ((~g28835));
assign g10085 = (g5556&g2483);
assign g10674 = (g3834&g5320);
assign g11877 = ((~g11111));
assign g14963 = ((~II21364));
assign g28848 = (g27875&g28610);
assign g12966 = (g7926&g10189);
assign g27425 = (g18025&g27138);
assign g16438 = (g2594&g12122);
assign g6103 = ((~II14624));
assign g24330 = ((~II31664));
assign g12695 = ((~II19787));
assign g24633 = (g24094)|(g20842);
assign g14894 = (g3940&g13148);
assign g29311 = ((~II38466));
assign g30780 = ((~g30625)&(~g22387));
assign g22710 = ((~II29386));
assign g30069 = ((~g29822)&(~g29828));
assign g10952 = ((~II17849));
assign g4214 = ((~g164));
assign g8263 = ((~II15457));
assign g19401 = ((~II25826));
assign g19543 = ((~II25966));
assign II36237 = ((~g27662));
assign g28617 = ((~g27858));
assign g9047 = (g6448&g7616);
assign g29392 = ((~g29042));
assign g12211 = ((~g8403));
assign g10936 = ((~II17831));
assign g18035 = (g5089&g15625);
assign II37858 = ((~g28501));
assign g27293 = ((~g27027)&(~g26357));
assign g9581 = (g6519&g8212);
assign g5297 = ((~II13849));
assign g27152 = ((~g23467)&(~g26062));
assign g15781 = (g7971&g13330);
assign g9033 = (g6643&g567);
assign g26271 = (g25907&g9468);
assign g24266 = ((~II31472));
assign g24527 = ((~g15509)&(~g23878));
assign II23000 = ((~g13872))|((~II22998));
assign g25565 = (g24496&g20466);
assign g16035 = ((~g12752));
assign g27082 = (g22016&g26639);
assign II13242 = ((~g2879));
assign g8939 = (g7195&g1874);
assign g17854 = (g4836&g15499);
assign g26687 = ((~II34668));
assign II23181 = ((~g13942))|((~II23179));
assign II36588 = ((~g27293));
assign g30207 = ((~g30028));
assign g16284 = (g8304&g11920);
assign g15329 = ((~II21598));
assign g24363 = ((~II31763));
assign II20580 = ((~g13364));
assign g12866 = ((~g8459)&(~g8482)&(~g8497));
assign g28404 = (g7792&g27843);
assign II31571 = ((~g24051));
assign g18204 = (g5243&g15726);
assign II32528 = ((~g24078))|((~II32526));
assign II18794 = ((~g10973));
assign g22316 = ((~g21149));
assign II31250 = ((~g22953));
assign g27385 = ((~II35723));
assign g27270 = ((~g26998)&(~g26298));
assign g30346 = ((~II39863));
assign g17988 = ((~g14685));
assign g26677 = ((~g25238)&(~g10340));
assign g26388 = (g5000&g25691);
assign g29636 = ((~II39026));
assign II39160 = ((~g29620));
assign g26665 = ((~g25348)&(~g17143));
assign g23983 = ((~g4809)&(~g22990));
assign g24908 = (g7342&g23882);
assign g15788 = ((~g12657))|((~g6574));
assign g18332 = ((~II24339))|((~II24340));
assign g11815 = ((~g9622)&(~g9746)&(~g9868));
assign II38731 = ((~g29328));
assign II25939 = ((~g2156))|((~II25938));
assign II15787 = ((~g6000));
assign II29304 = ((~g20945));
assign g20739 = ((~II27328));
assign g7715 = ((~g1697));
assign g21564 = (g13886&g14153&g19799&II28096);
assign II20021 = (g9941&g9857&g9737&g9613);
assign g29797 = ((~II39243));
assign g5104 = ((~g2436));
assign g23247 = ((~II30194));
assign g11447 = ((~II18411));
assign g22680 = ((~g20858))|((~g20928));
assign g11205 = ((~II18127));
assign g12448 = ((~II19618));
assign g21429 = ((~II27976));
assign g7748 = ((~g2393));
assign g17387 = ((~II23475));
assign g5425 = ((~II13987));
assign g25038 = ((~g23803))|((~g5556));
assign II30914 = ((~g22125));
assign II33535 = ((~g24508));
assign g15685 = ((~II21936));
assign g26922 = ((~g26283));
assign II40856 = ((~g30739));
assign II16661 = ((~g3774));
assign II35900 = ((~g26786));
assign II32635 = ((~g23970))|((~II32633));
assign g23387 = ((~g18508))|((~g22852));
assign II16212 = ((~g5411));
assign g28154 = ((~g27401));
assign g9103 = (g3462&g7706);
assign II25846 = ((~g771))|((~g18358));
assign II29206 = ((~g20910));
assign II35283 = ((~g26031));
assign g23007 = ((~g21491));
assign II40853 = ((~g30732));
assign g19297 = (g18115)|(g18212);
assign g10614 = (g6945&g1303);
assign g28736 = ((~g28427)&(~g27913));
assign g10292 = (g6912&g4623);
assign g9226 = ((~g5434));
assign g16775 = ((~II22763));
assign g25112 = ((~g24043))|((~g2753));
assign g10209 = (g6713&g4509);
assign g29337 = (g29103&g29032);
assign g8871 = ((~II16131));
assign g16158 = (g5718&g11834);
assign II18365 = ((~g7391));
assign g25935 = ((~g25127)&(~g17031));
assign g13406 = ((~II20517));
assign II32880 = ((~g24581));
assign g27139 = ((~g26226));
assign g20990 = ((~g19803)&(~g17813));
assign g26585 = ((~g25593));
assign g21130 = ((~II27689));
assign g5335 = ((~g2522));
assign g26481 = ((~g25764));
assign g24958 = ((~g23478));
assign II21392 = ((~g13020));
assign g30450 = ((~II40008));
assign g15449 = ((~II21711));
assign II28491 = ((~g21327));
assign g30637 = ((~g16141)&(~g30410));
assign II19915 = ((~g8560));
assign II38885 = ((~g29192));
assign g27037 = ((~g24933)&(~g26028));
assign g15509 = (g5008&g13227);
assign g27447 = ((~g27066))|((~g5556));
assign g7924 = ((~g3048));
assign II30782 = ((~g22081));
assign g27026 = (g22009&g26595);
assign g9216 = ((~g5966));
assign II20685 = ((~g11671));
assign II27516 = ((~g20333));
assign g4376 = ((~g1113));
assign g26998 = (g23325&g26566);
assign II34692 = ((~g26102));
assign g19295 = ((~II25617))|((~II25618));
assign II18665 = ((~g8689));
assign II34957 = ((~g26541));
assign II17433 = ((~g3900));
assign g8251 = ((~II15433));
assign II39878 = ((~g30282));
assign g27580 = ((~g26878))|((~g744));
assign g13278 = ((~g10158));
assign g28959 = ((~II37928));
assign g21761 = ((~g20198))|((~g6519));
assign II28753 = ((~g21893))|((~g13541));
assign g15055 = ((~g11952));
assign g12780 = ((~g9187)&(~g9161));
assign II14541 = ((~g455));
assign g22585 = ((~II29151));
assign g29367 = ((~g28911));
assign g10862 = ((~II17715));
assign II33855 = ((~g25350));
assign g23890 = ((~II31152));
assign II23976 = ((~g14719));
assign g27370 = (g27126&g8874);
assign g26288 = (g4592&g25524);
assign g30405 = ((~g30008)&(~g30133));
assign g21634 = (g19084)|(g19534)|(g16560);
assign g8372 = ((~II15574));
assign g7922 = ((~II15238))|((~II15239));
assign g28314 = ((~II37191));
assign g21529 = ((~g19272));
assign g22648 = ((~II29262));
assign g26630 = ((~g25309)&(~g24585));
assign g24883 = ((~II32596))|((~II32597));
assign g11858 = ((~g11085));
assign II37942 = ((~g28501));
assign g8816 = (g7303&g8084);
assign g22703 = ((~II29369));
assign g23098 = ((~g21678));
assign II38677 = ((~g29400));
assign g10202 = (g6912&g4483);
assign II16315 = ((~g3774));
assign g13871 = (g7898&g12775);
assign g21096 = ((~g20013)&(~g20051)&(~g20087));
assign g21938 = (g5832&g20550);
assign g5972 = ((~g2195));
assign g29046 = ((~II38003));
assign II31721 = ((~g23601));
assign II17151 = ((~g7142))|((~II17149));
assign g30727 = ((~II40471));
assign g13213 = ((~g9749));
assign II26337 = ((~g16880));
assign g19619 = (g3981&g17372);
assign g10422 = (g3306&g4882);
assign g11674 = ((~g9676))|((~g3522));
assign g4911 = ((~II13677));
assign g16662 = ((~II22706))|((~II22707));
assign II16826 = (g5903&g4507&g4508&g5234);
assign II21884 = ((~g13136));
assign II32167 = ((~g24230));
assign II37415 = ((~g28179));
assign g12026 = ((~g10195)&(~g10280)&(~g10360));
assign g22812 = ((~II29600));
assign II19516 = ((~g10683));
assign g17974 = ((~g14001));
assign g29201 = ((~g15104)&(~g28910));
assign g19187 = (g18419)|(g17729);
assign g10728 = ((~g3866))|((~g7488));
assign g13067 = ((~g9968))|((~g7426));
assign g11395 = ((~II18353));
assign II17831 = ((~g7518));
assign g13262 = ((~g10087));
assign g8825 = ((~II16047));
assign g5802 = ((~g83));
assign II17012 = ((~g6751));
assign g4665 = ((~g1416));
assign g15477 = ((~II21736));
assign g27507 = ((~g26941)&(~g24657));
assign g9528 = ((~II16681));
assign II25792 = ((~g17954))|((~II25790));
assign g22043 = ((~g21310)&(~g19570));
assign g8955 = ((~II16261));
assign II15267 = ((~g1161));
assign g23228 = ((~II30137));
assign g12542 = ((~g8684));
assign II24157 = ((~g14322))|((~II24156));
assign II34438 = ((~g25936));
assign II36108 = ((~g27360));
assign g13180 = ((~g9401));
assign g25697 = (g7455&g25120);
assign g19112 = (g14657&g16633);
assign g30830 = ((~II40742));
assign g11748 = ((~g10901));
assign II40426 = ((~g30581));
assign g21392 = (g15118&g20387);
assign g20384 = ((~g17511));
assign g17307 = ((~II23395));
assign g17094 = ((~g15962)&(~g15942)&(~g15923));
assign g30016 = ((~g29531)&(~g29949));
assign g11379 = ((~II18335));
assign g9118 = (g7265&g7751);
assign g29087 = ((~g9488))|((~g28595));
assign g8369 = ((~II15571));
assign g8182 = ((~g3198));
assign g22954 = ((~g21739));
assign g10983 = ((~II17884));
assign II29129 = ((~g20753));
assign g21030 = ((~II27585));
assign g10390 = (g5512&g4824);
assign g12891 = ((~g8925));
assign II20505 = ((~g11264))|((~II20504));
assign g27030 = (g22083&g26601);
assign g27333 = ((~g27085)&(~g26447));
assign g30320 = ((~II39803));
assign II20394 = ((~g10331));
assign g30280 = ((~g16425)&(~g30114));
assign g20560 = ((~II27005));
assign g22916 = ((~g8296))|((~g21725));
assign g11129 = ((~II18043));
assign II21075 = ((~g12506));
assign II27727 = ((~g19070));
assign g4721 = ((~g2501));
assign g26910 = ((~II35109));
assign g10830 = ((~II17677));
assign g23510 = (g5890&g22753);
assign g24325 = ((~II31649));
assign g19737 = (g4363&g17582);
assign g5645 = ((~g101));
assign II15278 = ((~g2938))|((~II15276));
assign g29630 = ((~II39008));
assign II33282 = ((~g25096));
assign g30621 = ((~g30412)&(~g2608));
assign g12961 = ((~g9000));
assign g24302 = ((~II31580));
assign g19368 = ((~II25772))|((~II25773));
assign II18040 = ((~g7976));
assign g30856 = ((~II40820));
assign g11608 = ((~II18784));
assign g28437 = ((~II37386));
assign II31475 = ((~g23555));
assign g8482 = (g7085&g2300);
assign g15835 = ((~g12611))|((~g6519));
assign g19412 = ((~g16673));
assign II40438 = ((~g30583));
assign g13050 = ((~g9822))|((~g7230));
assign g26425 = (g25923&g9958);
assign g26069 = (g25949&g21130);
assign g25963 = (g24756&g11944);
assign g26745 = ((~II34842));
assign g12192 = ((~g10423)&(~g10485)&(~g10548));
assign g28987 = ((~g28666)&(~g13390));
assign g26688 = ((~II34671));
assign g14016 = ((~g12852));
assign g8258 = ((~II15442));
assign g4052 = ((~g1412));
assign g19247 = ((~II25506));
assign g29748 = ((~g6104)&(~g29583)&(~g25363));
assign g24518 = ((~II32042));
assign g13082 = (II20131&II20132);
assign g4073 = ((~g2220));
assign II30062 = ((~g22590));
assign II37467 = ((~g27760));
assign g7788 = ((~g1345));
assign g25991 = ((~II33825));
assign II34469 = ((~g25210));
assign g29289 = (g29030&g28883);
assign g5123 = ((~g2784));
assign g5789 = ((~g1886));
assign g26205 = ((~II34121));
assign g6517 = ((~g283));
assign g23584 = (g6167&g22470);
assign g10271 = (g7426&g4584);
assign g19520 = (g16974&g15003&g14936);
assign g8771 = ((~II15967));
assign II13652 = ((~g2170));
assign II18704 = ((~g11055));
assign g22687 = ((~g21926)&(~g19010));
assign g19635 = (g1319&g18811);
assign g10073 = (g7358&g4286);
assign g19173 = ((~g17636)&(~g15389));
assign g27694 = ((~II36093));
assign II16736 = (g5713&g5958&g4735&g4736);
assign g27148 = ((~g26393));
assign g27286 = ((~g27020)&(~g26340));
assign II17939 = ((~g6232));
assign g18424 = ((~II24444))|((~II24445));
assign g29813 = (g29760&g13869);
assign II19836 = ((~g8726));
assign g18179 = ((~g14153));
assign g10680 = (g6980&g5330);
assign g5902 = ((~g945));
assign g4092 = ((~g3074));
assign g11318 = ((~II18268));
assign g21042 = ((~g19882)&(~g15634));
assign II31616 = ((~g23619));
assign II35796 = ((~g27122));
assign g21082 = ((~g19941)&(~g18330));
assign g22400 = ((~g21235))|((~g14618))|((~g10754));
assign g30114 = (g29865&g11447);
assign g17186 = ((~g7949)&(~g14144));
assign g13636 = (g6205&g12493);
assign II16493 = ((~g7936));
assign II33798 = ((~g25109));
assign g21671 = ((~II28201));
assign g5126 = ((~g2789));
assign g28423 = (g17724&g28152);
assign II14783 = ((~g1520));
assign II33891 = ((~g25850));
assign gbuf45 = (g382);
assign II40895 = ((~g30826));
assign II39279 = ((~g29708));
assign II24279 = ((~g6284))|((~II24278));
assign g13087 = ((~g9534))|((~g6678));
assign g30085 = (g29829&g11092);
assign g29224 = ((~g28970)&(~g28481));
assign g9077 = (g6448&g7649);
assign g8601 = (g6643&g7153);
assign g12555 = ((~II19727));
assign g21351 = (g9174&g20349);
assign II24973 = ((~g15003));
assign g28648 = ((~g27965));
assign g21047 = ((~g19888)&(~g15651));
assign g4325 = ((~g36));
assign g11987 = ((~g10120)&(~g10209)&(~g10295));
assign g23969 = ((~g22852))|((~g13974));
assign g5896 = ((~g261));
assign g30679 = ((~g16429)&(~g30504));
assign II32490 = ((~g18131))|((~g24067));
assign II26682 = (g15003&g18796&g13774);
assign g19949 = (g5293&g18278);
assign g20662 = ((~II27253));
assign g20597 = ((~II27116));
assign g22662 = ((~II29288));
assign g29693 = ((~II39133));
assign g29626 = (g29318&g11478);
assign II20538 = ((~g13384));
assign g19641 = ((~g16943));
assign g5153 = ((~g1136));
assign II34767 = ((~g26246));
assign II15237 = ((~g2963))|((~g2966));
assign g5679 = ((~g506));
assign g12654 = ((~II19774));
assign II36797 = ((~g27346));
assign II14885 = ((~g1786));
assign g6711 = ((~g281));
assign g22911 = ((~g21246))|((~g771));
assign g26391 = (g25923&g9876);
assign II18079 = ((~g6783));
assign g12849 = ((~g8433)&(~g8464)&(~g8485));
assign g12382 = ((~II19542));
assign g23904 = (g3010&g22750);
assign g24830 = ((~II32423))|((~II32424));
assign g27130 = ((~g26451))|((~g5556));
assign g27160 = ((~g23476)&(~g26069));
assign II31730 = ((~g23627));
assign II21432 = ((~g13044));
assign II22963 = ((~g9161))|((~II22962));
assign g23688 = (g23106)|(g21906);
assign g17528 = (g4257&g15201);
assign g13448 = ((~II20643));
assign II21267 = ((~g11663));
assign g13106 = ((~g9822))|((~g7358));
assign g5176 = ((~g1958));
assign g28419 = ((~g28151));
assign g21358 = ((~II27897));
assign g5834 = ((~g2175));
assign II24374 = ((~g9310))|((~II24372));
assign g18070 = ((~g15854));
assign g27103 = (g5235&g26461);
assign gbuf38 = (g350);
assign g28464 = (g26121&g28169);
assign II16012 = ((~g5390));
assign II29162 = ((~g20897));
assign g14008 = ((~II21037));
assign g23661 = ((~II30797));
assign g30907 = ((~II40973));
assign g25251 = ((~g24824)&(~g23679));
assign II15605 = ((~g6574));
assign g27886 = ((~g27632)&(~g24627));
assign g20331 = ((~g17357));
assign g10435 = (g3366&g4899);
assign II15559 = ((~g7015));
assign II23124 = ((~g9374))|((~II23123));
assign II21601 = ((~g13087));
assign g4243 = ((~g851));
assign g29513 = ((~II38869));
assign II38743 = ((~g29267));
assign II23094 = ((~g9326))|((~II23093));
assign g8458 = (g7085&g2291);
assign g21449 = ((~II27992));
assign g16852 = ((~II22828));
assign g28283 = ((~II37098));
assign g5658 = (g1012&g1036);
assign II18408 = ((~g6574));
assign g13365 = (g5785&g11389);
assign g26596 = ((~g13853)&(~g25304));
assign II18073 = ((~g6945));
assign II27011 = ((~g19546));
assign g24029 = (g2900&g22903);
assign II29010 = ((~g21724));
assign g26955 = (g6157&g26533);
assign g15731 = ((~II21979));
assign g9711 = ((~g5735));
assign g18605 = ((~II24703))|((~II24704));
assign II28031 = ((~g19172));
assign g22075 = ((~g21339)&(~g19618));
assign II38647 = ((~g29306));
assign g7900 = ((~g3075));
assign II21705 = ((~g11700));
assign gbuf40 = (g357);
assign g10443 = (g6751&g4925);
assign g10904 = ((~g5922));
assign II32857 = ((~g23748));
assign g20613 = ((~II27164));
assign II22926 = ((~g14091))|((~II22924));
assign II28217 = ((~g14194))|((~g19471));
assign g24409 = ((~II31901));
assign II30676 = ((~g22048));
assign g28027 = (g27590&g9895);
assign g12882 = ((~g8921));
assign II34135 = ((~g25229));
assign II22771 = ((~g14677));
assign II22539 = ((~g14882));
assign g23694 = ((~II30864));
assign g13129 = ((~g9822))|((~g7230));
assign gbuf29 = (g452);
assign g28432 = ((~II37379));
assign g22218 = ((~g21639)&(~g19949));
assign II23851 = ((~g15930));
assign II24195 = ((~g13927))|((~II24194));
assign II40300 = ((~g30485));
assign g21659 = ((~g20164))|((~g6314));
assign g4728 = ((~g2780));
assign g9757 = ((~g5601));
assign g13918 = ((~g11830));
assign g29790 = (g29491&g10918);
assign g25479 = ((~II33307));
assign g15738 = ((~g12415));
assign II38505 = ((~g28774));
assign g30808 = ((~II40676));
assign g20874 = ((~g17301)&(~g19594));
assign g18311 = (g5306&g15766);
assign g29767 = ((~g29468)&(~g19143));
assign g12170 = ((~g10395)&(~g10458)&(~g10520));
assign g28525 = ((~g27245)&(~g27726));
assign g24575 = ((~g23972)&(~g22874));
assign g15959 = ((~g2814)&(~g13082));
assign g27171 = ((~II35376));
assign g8200 = ((~g168));
assign g19702 = (g4237&g17514);
assign g26662 = ((~g25877));
assign g28322 = (g27937&g13868);
assign gbuf22 = (g138);
assign II35431 = ((~g26868));
assign g10360 = (g3306&g4737);
assign g23279 = ((~II30290));
assign g4121 = ((~g705));
assign g30944 = (g30935&g20666);
assign g19809 = (g1352&g18898);
assign g5469 = ((~g3085));
assign g11889 = ((~g9887)&(~g10007)&(~g10101));
assign g28071 = ((~II36656));
assign II23383 = ((~g15811));
assign g17402 = ((~II23490));
assign II31008 = ((~g22150));
assign g28104 = (g27608&g10232);
assign g19804 = (g679&g18893);
assign g7629 = ((~g403));
assign g14062 = ((~g12880));
assign g21022 = ((~g19854)&(~g15572));
assign II35172 = ((~g26272));
assign II40537 = ((~g30694));
assign g8099 = ((~g3061));
assign II39475 = ((~g29938));
assign g16865 = (g6896&g14881);
assign g5761 = ((~g797));
assign II18386 = ((~g3254));
assign g16988 = (g7842&g15261);
assign g5720 = ((~g986));
assign II18644 = ((~g8937));
assign g28392 = ((~g27886)&(~g22344));
assign II25572 = ((~g740))|((~II25571));
assign g27502 = ((~II35856));
assign g13674 = (g6431&g12530);
assign g8553 = (g6574&g1585);
assign g18945 = ((~g15667));
assign g14881 = ((~g11923));
assign g20313 = ((~g17310));
assign g26220 = ((~II34150));
assign g17247 = ((~g16050)&(~g16070));
assign g30698 = (g30383&g11126);
assign II18061 = ((~g3410));
assign g22151 = ((~g21421)&(~g19747));
assign g14165 = ((~g11975));
assign g6369 = ((~II14742));
assign g23729 = ((~II30911));
assign g30372 = (g8594&g30228);
assign g28376 = (g744&g27990);
assign g22166 = ((~g21445)&(~g19779));
assign II29026 = ((~g21737));
assign g26982 = (g21983&g26556);
assign g29424 = ((~II38653));
assign II19820 = ((~g10560));
assign g13170 = ((~g9323));
assign g28725 = ((~g28499));
assign g21002 = ((~g19819)&(~g15505));
assign g21875 = ((~g18531))|((~g19235))|((~g19245));
assign g18856 = ((~g15340));
assign g5401 = ((~II13919));
assign g13862 = (g5366&g12743);
assign II19315 = ((~g10424));
assign g6978 = ((~g1245));
assign g19158 = ((~II25355));
assign g21079 = ((~g20550));
assign g26823 = ((~g15437)&(~g26353));
assign g18504 = ((~II24554))|((~II24555));
assign II16650 = ((~g3618));
assign II37760 = ((~g28540));
assign g12790 = ((~g8847));
assign g23919 = (g22666)|(g23140);
assign g15550 = ((~II21806));
assign II34369 = ((~g25263));
assign g28062 = ((~II36633));
assign g29466 = (g8587&g29265);
assign g19233 = (g18302)|(g18383);
assign g10901 = ((~II17774));
assign II25811 = ((~g17993))|((~II25809));
assign g15196 = (g4375&g13178);
assign g15923 = ((~g11630));
assign g12426 = ((~II19576));
assign g17566 = ((~g16346));
assign g13568 = ((~g11627));
assign g14442 = ((~g11768));
assign g28762 = ((~g28446)&(~g27938));
assign g10389 = (g7015&g4821);
assign g20156 = (g16809&g3185);
assign g17142 = ((~II23162))|((~II23163));
assign g29487 = (g21580&g29292);
assign II14819 = ((~g1092));
assign g28584 = (g27756)|(g25874);
assign g16177 = ((~g12895));
assign g28005 = ((~II36496));
assign g7812 = ((~g2398));
assign g7827 = ((~g478));
assign II35879 = ((~g26814));
assign II29191 = ((~g20901));
assign g19021 = ((~II25126));
assign g11498 = ((~II18470));
assign g30248 = ((~g16139)&(~g30081));
assign g16040 = ((~g12759));
assign II25399 = ((~g18794));
assign g24648 = ((~g23470));
assign g11717 = ((~g9676))|((~g3522));
assign g24335 = ((~II31679));
assign g29433 = ((~II38680));
assign g19595 = ((~II26025));
assign II20425 = ((~g10842));
assign g26604 = ((~g25658));
assign g22832 = ((~II29619));
assign g12950 = ((~g8990));
assign g27823 = ((~g27632)&(~g1216));
assign II20117 = ((~g10876));
assign g26883 = ((~II35076));
assign g23242 = ((~II30179));
assign g10047 = (g6713&g1107);
assign g9507 = ((~g5953));
assign g12264 = ((~g8449));
assign II15584 = ((~g3254));
assign g6943 = ((~g801));
assign g20438 = ((~g17710));
assign g26426 = (g5115&g25755);
assign II36502 = ((~g27269));
assign II36891 = ((~g28004));
assign g26446 = (g5179&g25790);
assign g8027 = ((~g3069));
assign g17240 = ((~II23326));
assign g19151 = ((~II25344));
assign g9050 = ((~g5731));
assign II23521 = ((~g13518));
assign II22836 = ((~g13571));
assign g24820 = ((~II32401))|((~II32402));
assign g19838 = ((~II26276));
assign g20360 = ((~II26777));
assign g27514 = ((~II35876));
assign g19093 = (g17218&g16572);
assign g28353 = ((~g15666)&(~g28073));
assign g9425 = ((~g5346));
assign g23050 = ((~II29797));
assign g13699 = ((~g13252));
assign g26884 = ((~II35079));
assign g29769 = ((~g29470)&(~g19148));
assign g4753 = ((~g599));
assign g19864 = (g18247&g16131);
assign II30152 = ((~g22713));
assign g27533 = ((~II35915));
assign g12177 = ((~g8375));
assign II40456 = ((~g30668));
assign g18622 = ((~g14613));
assign g7822 = ((~g510));
assign II26541 = (g18538&g18484&g18406);
assign g19494 = ((~g18218));
assign g16415 = (g5956&g12077);
assign g19279 = (g17942)|(g18030);
assign g27703 = ((~II36120));
assign g19742 = (g1332&g18857);
assign g12822 = ((~II19883));
assign g13859 = ((~g11608));
assign g30363 = ((~II39902));
assign g24067 = ((~g22887))|((~g14486));
assign g8083 = ((~g1862));
assign g30354 = ((~II39881));
assign g29475 = (g21544&g29272);
assign g29972 = ((~II39454));
assign II30050 = ((~g22619));
assign g3410 = ((~II13179));
assign II39133 = ((~g29609));
assign g11566 = ((~II18674));
assign g24486 = ((~g23643)&(~g22577));
assign g24056 = ((~g22887))|((~g14554));
assign g10185 = ((~II17150))|((~II17151));
assign g15337 = (g4650&g13198);
assign II29562 = ((~g21035));
assign g25033 = ((~g23955))|((~g6751));
assign g19929 = (g2753&g18965);
assign II37897 = ((~g28501));
assign g15525 = ((~g12336));
assign g24586 = ((~II32150));
assign g13511 = ((~g12611))|((~g3410));
assign g26192 = ((~II34102));
assign g24492 = ((~g23689)&(~g22610));
assign g28253 = ((~II37008));
assign g6220 = ((~g2598));
assign g30125 = ((~II39638));
assign g25968 = (g24871&g11986);
assign gbuf182 = (g2363);
assign g23216 = ((~II30101));
assign g24520 = ((~g23829)&(~g22707));
assign g28399 = (g7776&g27820);
assign g13962 = ((~g11864));
assign g25059 = ((~g23984))|((~g7195));
assign g28729 = (g28606&g16794);
assign g26504 = (g5338&g25877);
assign g21203 = (g20178&g12409);
assign g15126 = (g4249&g13169);
assign II33861 = ((~g25744));
assign II17948 = ((~g6643));
assign g12596 = ((~g8748));
assign II25607 = ((~g17825))|((~II25605));
assign g11675 = ((~g9107)&(~g9114)&(~g9120));
assign II36090 = ((~g27502));
assign g20410 = ((~g17604));
assign g27797 = ((~II36246));
assign g26891 = ((~g25561)&(~g26345));
assign g11824 = ((~g11022));
assign II21108 = ((~g13150));
assign g24857 = ((~II32510))|((~II32511));
assign g26489 = ((~II34453));
assign g7760 = ((~g2392));
assign g12220 = ((~g8418));
assign g21308 = (g9374&g20303);
assign g21483 = ((~II28019));
assign g4587 = ((~g2799));
assign g25395 = ((~g24916));
assign g9260 = ((~II16514));
assign II28981 = ((~g21667));
assign g30467 = (g30179&g11274);
assign g16065 = ((~g12811));
assign II23599 = ((~g15887));
assign g6284 = ((~g640));
assign II15568 = ((~g3722));
assign II23490 = ((~g15823));
assign g9884 = ((~g6310));
assign g12457 = ((~g9009)&(~g9033)&(~g9048));
assign g16412 = ((~g12565))|((~g3254));
assign g13159 = ((~g9245));
assign II40754 = ((~g30666));
assign g13756 = ((~g12448));
assign g24448 = ((~g23923))|((~g3338));
assign g26125 = ((~II34020));
assign g26348 = (g4829&g25615);
assign g15792 = ((~g12426));
assign g19253 = (g17121)|(g17085)|(II25516);
assign g26020 = ((~II33912));
assign g14408 = ((~g12112));
assign II40742 = ((~g30662));
assign g15248 = ((~II21531));
assign g27632 = ((~II36032));
assign g19269 = (g17049)|(g17020)|(II25554);
assign g19193 = (g18492)|(g17998);
assign II28512 = ((~g21496));
assign g20810 = ((~II27399));
assign g9504 = ((~g6149));
assign g4620 = ((~g728));
assign g12218 = ((~g8411));
assign g29917 = ((~II39348))|((~II39349));
assign g19760 = (g2727&g18864);
assign g30762 = (g30608&g20830);
assign g21168 = ((~g20162)&(~g20191)&(~g20220));
assign II21666 = ((~g13100));
assign g15698 = ((~g12389));
assign g27253 = ((~g26965)&(~g26212));
assign g26989 = ((~g26663)&(~g21913));
assign II22584 = ((~g15989));
assign g10282 = (g3306&g444);
assign g30266 = ((~g16359)&(~g30100));
assign g10119 = (g6519&g4369);
assign g11832 = ((~g9662)&(~g9777)&(~g9905));
assign g16429 = (g5973&g12115);
assign g26150 = ((~II34044));
assign g23274 = ((~II30275));
assign g24471 = ((~g23803))|((~g3774));
assign gbuf178 = (g2355);
assign g22387 = ((~g21250));
assign g13295 = (g1679&g11170);
assign g21892 = (g19288&g13011);
assign g24236 = (g22243&g11157);
assign g18963 = ((~g15734));
assign g8062 = ((~g169));
assign g30100 = (g29865&g11306);
assign g15729 = (g5304&g13297);
assign g26873 = ((~g25483)&(~g26260));
assign g13044 = ((~g9534))|((~g6678));
assign g20980 = ((~g19787)&(~g15435));
assign g22228 = (g21716&g12136);
assign II34641 = ((~g26086));
assign g16475 = ((~II22527));
assign II32949 = ((~g24605));
assign g10835 = ((~g5788)&(~g5827)&(~g5872));
assign g19881 = (g2059&g18935);
assign g20687 = ((~II27278));
assign II14295 = ((~g3228));
assign g15343 = ((~II21612));
assign g29670 = ((~g29529)&(~g29302));
assign g10637 = (g3806&g5269);
assign g30454 = (g30147&g11199);
assign g30672 = ((~g16401)&(~g30489));
assign II40763 = ((~g30729));
assign g16659 = ((~II22702));
assign g28670 = (g27798&g21935);
assign g26974 = (g26157)|(g23147);
assign g27770 = (g5642&g27449);
assign g12166 = ((~II19345));
assign g13990 = ((~g8594))|((~g12495));
assign g19260 = (g16749&g3124);
assign g27542 = ((~II35930));
assign g15813 = ((~g13011));
assign g29290 = ((~g28814));
assign g16223 = ((~g12006));
assign g22029 = ((~g21292)&(~g19555));
assign g19652 = ((~II26078));
assign g19822 = (g4708&g17779);
assign g8687 = (g3338&g7827);
assign g21444 = (g6568&g20427);
assign g29157 = ((~II38214));
assign g17544 = (g4292&g15231);
assign II35762 = ((~g26918));
assign g16419 = (g5960&g12085);
assign II20295 = ((~g10015));
assign g25088 = ((~g23950))|((~g679));
assign II27122 = ((~g19595));
assign g26543 = ((~g25476));
assign g5024 = ((~g449));
assign II16514 = ((~g5473));
assign g25524 = ((~II33352));
assign g21266 = ((~g20040));
assign g16075 = ((~g11861));
assign g7892 = ((~g2553));
assign II21739 = ((~g13091));
assign g25130 = ((~II32868));
assign g20316 = ((~g17318));
assign g28686 = ((~II37605));
assign II33437 = ((~g25046));
assign g23065 = ((~II29812));
assign g3951 = ((~g840));
assign II36397 = ((~g27574));
assign II15810 = ((~g3338));
assign g29910 = (g29779&g9961);
assign g30650 = ((~g16264)&(~g30451));
assign g8447 = (g6783&g1606);
assign g21445 = (g9795&g20428);
assign g21968 = ((~g21234)&(~g19476));
assign g21267 = (g20318&g16764&g16708);
assign g25672 = ((~II33498));
assign g18240 = ((~g14606)&(~g16094));
assign II20616 = ((~g13294));
assign g19217 = ((~II25456));
assign II23095 = ((~g13935))|((~II23093));
assign g30657 = ((~g16311)&(~g30461));
assign g24459 = ((~g23955))|((~g3494));
assign g8191 = ((~g147));
assign g19038 = ((~II25177));
assign II31892 = ((~g23801));
assign g28268 = ((~II37053));
assign II33912 = ((~g25891));
assign II24252 = ((~g7329))|((~II24251));
assign g19757 = (g4427&g17627);
assign II37746 = ((~g28595));
assign g30683 = ((~g16453)&(~g30334));
assign gbuf105 = (g1256);
assign g28189 = ((~g27359)&(~g26853));
assign g30077 = (g29823&g10963);
assign g27118 = ((~g26320))|((~g5438));
assign g20019 = (g17830)|(g18492)|(II26461);
assign g24450 = ((~g23748))|((~g3618));
assign II32085 = ((~g24179));
assign g29268 = ((~g28751));
assign g15780 = (g7471&g3032&II22028);
assign g19186 = (g18419)|(g17887);
assign g11673 = ((~g9676))|((~g3522));
assign II20355 = ((~g10229));
assign g20198 = ((~II26642));
assign II29954 = ((~g22611));
assign II21962 = ((~g13004));
assign II31559 = ((~g24233));
assign g28009 = (g14454&g27510);
assign g24090 = ((~g22887))|((~g14217));
assign II31469 = ((~g23546));
assign g9569 = ((~g5683));
assign gbuf93 = (g1067);
assign g20995 = ((~g19809)&(~g17837));
assign g29897 = ((~g29686));
assign g5729 = (g1018&g1053);
assign g15326 = ((~II21595));
assign II17184 = ((~g3494));
assign gbuf117 = (g1206);
assign g17324 = ((~II23412));
assign II18396 = ((~g3410));
assign g28634 = ((~g28185)&(~g17001));
assign g23687 = (g22668&g17570);
assign g24760 = (g9427&g24112);
assign g28243 = ((~II36978));
assign II37851 = ((~g28668));
assign g12441 = ((~g8594)&(~g10767));
assign II14163 = ((~g113));
assign g27766 = ((~g27554)&(~g27104));
assign g16277 = (g5634&g13275);
assign g7911 = ((~II15230));
assign g14507 = ((~g12179));
assign g6201 = ((~g646));
assign g5925 = ((~g189));
assign II27832 = ((~g19921));
assign II21326 = ((~g12378));
assign g26400 = (g5041&g25711);
assign II31844 = ((~g23633));
assign g30017 = ((~g29532)&(~g29950));
assign g10585 = (g3678&g5187);
assign g11092 = ((~II18004));
assign g11879 = ((~g11117));
assign g11845 = ((~II19025));
assign g29010 = ((~II37973));
assign g26373 = (g4925&g25664);
assign g13815 = (g7139&g12560);
assign II27246 = ((~g19335));
assign g15787 = ((~g12611))|((~g6519));
assign g15641 = ((~II21894));
assign g20894 = ((~g19629)&(~g17450));
assign g18821 = ((~g13740)&(~g11926));
assign g27497 = ((~II35849));
assign g4623 = ((~g733));
assign g19251 = ((~g16540));
assign II25635 = ((~g17640))|((~II25633));
assign II36315 = ((~g27575))|((~II36314));
assign g5680 = ((~g749));
assign g4197 = ((~g2251));
assign II32617 = ((~g24091))|((~II32615));
assign g13825 = ((~g12462));
assign g12993 = ((~g9035));
assign g3554 = ((~II13197));
assign g15842 = ((~g13332))|((~g12392));
assign g8892 = (g3338&g496);
assign II37311 = ((~g27897))|((~g27883));
assign g23251 = ((~II30206));
assign II13207 = ((~g1782));
assign g24815 = ((~g23448));
assign g4009 = ((~g174));
assign g3366 = ((~II13173));
assign g24264 = ((~II31466));
assign g18941 = ((~g15652));
assign g16360 = ((~g13063));
assign II19898 = ((~g10664));
assign g10174 = (g5556&g2492);
assign II18308 = ((~g6448));
assign g12242 = ((~II19415));
assign g29582 = ((~g29409)&(~g17100));
assign g29107 = ((~g9941))|((~g28595));
assign g28372 = ((~II37273));
assign g5765 = ((~g797));
assign g18830 = ((~g15225));
assign g27526 = ((~II35900));
assign g15811 = ((~g12711))|((~g6838));
assign g5874 = ((~g1888));
assign gbuf75 = (g963);
assign g21189 = ((~g20098)&(~g20061));
assign g15106 = ((~II21426));
assign g19248 = (g16662&g8817);
assign g24222 = ((~g17017)&(~g22272));
assign g28396 = (g7754&g27806);
assign g14669 = ((~II21256));
assign g20293 = (g14922&g18765&g13724&g16360);
assign g11681 = ((~g9111)&(~g9118)&(~g9123));
assign g20973 = ((~g19775)&(~g17753));
assign g4956 = ((~g1957));
assign gbuf179 = (g2357);
assign II21758 = ((~g13094));
assign II21297 = ((~g11687));
assign g24791 = ((~II32334))|((~II32335));
assign g14297 = (g7757&g12993);
assign II26266 = ((~g17791));
assign g28694 = ((~II37629));
assign g17022 = (g7892&g15439);
assign g29982 = (g29893&g8336);
assign II27976 = ((~g19957));
assign g27383 = ((~g27133));
assign g23348 = ((~g22195)&(~g10340));
assign II33312 = ((~g25014));
assign II31760 = ((~g23713));
assign II34266 = ((~g25255));
assign g29834 = (g29713&g22366);
assign g8780 = ((~II15978));
assign II31796 = ((~g23508));
assign g22148 = ((~g21414)&(~g19739));
assign g30520 = ((~II40140));
assign g30513 = ((~II40119));
assign g21750 = ((~g20255))|((~g7085));
assign g18401 = ((~g16233)&(~g7134));
assign g26438 = (g5159&g25776);
assign g13032 = (g3996&g10545);
assign II37173 = ((~g28132));
assign g4091 = ((~g2864));
assign II36679 = ((~g27316));
assign g12065 = ((~g11401));
assign g5983 = ((~g879));
assign g29817 = (g29709&g20694);
assign II19513 = ((~g10664));
assign II32281 = ((~g23950));
assign g13884 = (g7594&g12807);
assign g13294 = ((~II20355));
assign g11942 = ((~g11219));
assign g19166 = (g17212&g8637);
assign g7194 = ((~II14925));
assign II22936 = ((~g9150))|((~g13906));
assign II27614 = ((~g20067));
assign II33834 = ((~g25667));
assign g13526 = ((~g12711))|((~g3722));
assign II15205 = ((~g2969))|((~II15204));
assign g10681 = (g3650&g2000);
assign g6837 = ((~II14839));
assign g21276 = (g20337&g16791&g16739);
assign II25605 = ((~g744))|((~g17825));
assign g20134 = (g18337&g9506);
assign g20601 = ((~II27128));
assign II29226 = ((~g20917));
assign II31652 = ((~g23784));
assign g8075 = ((~g1547));
assign II19816 = ((~g10703));
assign g24338 = ((~II31688));
assign g14061 = ((~g11928));
assign II20679 = ((~g11641));
assign g25923 = ((~g24963));
assign II26420 = ((~g17042));
assign g13126 = ((~g9676))|((~g7162));
assign g25149 = ((~II32925));
assign g29495 = ((~II38801));
assign g24776 = (g9507&g24129);
assign g11722 = ((~g9676))|((~g3522));
assign g10784 = ((~g5630)&(~g5649)&(~g5676));
assign g30583 = ((~II40303));
assign g30699 = ((~g13914)&(~g30387));
assign g25004 = ((~g23644))|((~g6448));
assign g13248 = ((~II20299));
assign g6942 = ((~g279));
assign g30730 = ((~II40478));
assign II18770 = ((~g10333));
assign g19199 = ((~II25432));
assign g28784 = ((~g28468)&(~g27970));
assign g9767 = ((~II16811));
assign g23306 = ((~II30371));
assign g27999 = ((~II36486));
assign g23088 = ((~g21655));
assign g8385 = (g3254&g228);
assign II25654 = ((~g1430))|((~II25653));
assign II16641 = ((~g6713));
assign II23314 = ((~g15720));
assign II30888 = ((~g22115));
assign g26769 = (g14753&g26525);
assign g17619 = (g4415&g15290);
assign g26999 = (g21983&g26567);
assign II24646 = ((~g14385))|((~g9795));
assign g21882 = ((~g13862)&(~g19248));
assign g23453 = ((~II30483));
assign g12216 = ((~g10462)&(~g10523)&(~g10585));
assign g16130 = ((~g12868));
assign g4526 = ((~g1415));
assign g7158 = ((~g1171));
assign g8757 = ((~II15949));
assign g30062 = ((~g29810)&(~g29815));
assign g30007 = (g29905&g8494);
assign g12196 = ((~g8388));
assign g22551 = ((~II29107));
assign g16238 = (g12275&g11066);
assign g21285 = ((~II27832));
assign II23358 = ((~g16442));
assign g22833 = ((~II29622));
assign g26849 = ((~II35000));
assign II16267 = ((~g5473));
assign II22964 = ((~g13885))|((~II22962));
assign g11595 = ((~II18761));
assign II29588 = ((~g21046));
assign II20031 = ((~g10003))|((~g9883));
assign g25648 = ((~g24720)&(~g24500));
assign II16578 = ((~g6448));
assign II34845 = ((~g26496));
assign g28128 = ((~g27528));
assign g18638 = (g13805&g13840&II24758);
assign g4644 = ((~g1045));
assign g28354 = ((~g15670)&(~g28079));
assign g19857 = (g4854&g17859);
assign II35667 = ((~g27120));
assign II15475 = ((~g3246));
assign g13724 = ((~g12470));
assign g28471 = (g18190&g27956);
assign g24099 = ((~g22412));
assign g23195 = ((~II30038));
assign g23795 = (g18110&g23028);
assign II24612 = ((~g15814))|((~II24611));
assign II19274 = ((~g10560));
assign II38477 = ((~g28760));
assign g25023 = ((~g23955))|((~g6945));
assign g25066 = ((~g23984))|((~g7195));
assign g14412 = ((~g12113));
assign g11514 = ((~II18518));
assign II13200 = ((~g1547));
assign II14665 = ((~g3147));
assign g25180 = ((~II33016));
assign II26621 = (g14863&g18735&g18789);
assign g15826 = ((~g12711))|((~g6838));
assign g26000 = ((~II33852));
assign g4839 = ((~g2094));
assign g18448 = ((~g13974));
assign g18030 = ((~II24062))|((~II24063));
assign g4208 = ((~g133));
assign g20517 = ((~g18450));
assign g26534 = ((~g25321)&(~g8869));
assign II22560 = ((~g14796));
assign g13076 = ((~g10818));
assign g22434 = ((~II28978));
assign II32895 = ((~g24816));
assign g26621 = ((~g25711));
assign g25365 = (g24700&g18236);
assign II19767 = ((~g8726));
assign g21031 = ((~g19869)&(~g17989));
assign g7936 = ((~II15256));
assign II25681 = ((~g70))|((~g17974));
assign g20676 = ((~II27267));
assign g21057 = ((~II27614));
assign g16636 = ((~II22679));
assign g17557 = ((~II23645));
assign g19078 = ((~g18619));
assign II31643 = ((~g23737));
assign g11507 = ((~II18497));
assign g26752 = ((~II34863));
assign II28458 = ((~g20971));
assign g28017 = ((~II36524));
assign g10606 = ((~g8074));
assign g22013 = ((~g21277)&(~g19548)&(~g19551));
assign g20054 = ((~g19001)&(~g16867));
assign g29521 = (g28733&g29362);
assign g18585 = ((~g14135));
assign g28086 = (g27608&g10158);
assign g17508 = (g4225&g15179);
assign g12534 = ((~II19702));
assign g19387 = ((~g16567));
assign g13355 = (g5756&g11355);
assign g19080 = (g18708&g14991&g13724&g16313);
assign g16471 = ((~II22515));
assign II39341 = ((~g29741))|((~II39339));
assign g28103 = ((~II36744));
assign g27094 = ((~g4809)&(~g26090));
assign g20628 = ((~II27209));
assign II14650 = ((~g525));
assign II24091 = ((~g13886))|((~g15096));
assign g20312 = ((~g17307));
assign g21258 = ((~g20002));
assign II33355 = ((~g25012));
assign II32175 = ((~g24235));
assign g14650 = ((~II21249));
assign g5141 = ((~II13775));
assign g22880 = ((~g19468))|((~g20904));
assign g18142 = ((~g14124));
assign II25673 = ((~g18469))|((~II25671));
assign g14206 = ((~g11993));
assign g30044 = ((~g29916));
assign g16123 = ((~g12923))|((~g1319));
assign II40685 = ((~g30643));
assign g5269 = ((~g2652));
assign g16862 = ((~II22842));
assign g8766 = ((~II15958));
assign g6065 = ((~II14574));
assign g21957 = ((~II28497));
assign II24487 = ((~g9391))|((~II24485));
assign g22291 = (g21766&g12318);
assign II23611 = ((~g14966));
assign II29119 = ((~g20883));
assign gbuf46 = (g387);
assign g28320 = (g27854&g20637);
assign g28527 = ((~II37474));
assign g20327 = ((~g17342));
assign II16782 = ((~g6083));
assign g26628 = ((~g25738));
assign g14493 = ((~II21208));
assign g15505 = (g4842&g12830);
assign g11993 = ((~g10153)&(~g10224)&(~g10310));
assign g30960 = ((~g30924)&(~g30950));
assign II25723 = ((~g18341))|((~II25721));
assign II14553 = ((~g1056));
assign g12290 = ((~g10573)&(~g10616)&(~g10652));
assign g10963 = ((~II17854));
assign g7539 = ((~g2528));
assign II18353 = ((~g3722));
assign g30927 = ((~II41018))|((~II41019));
assign g4603 = ((~g577));
assign II41102 = ((~g30969));
assign II40558 = ((~g30605))|((~g30597));
assign g26392 = (g5005&g25694);
assign II36792 = ((~g27345));
assign g30839 = ((~II40769));
assign g15488 = ((~II21747));
assign g27162 = ((~g26461));
assign II29277 = ((~g20935));
assign g30853 = ((~II40811));
assign II16050 = ((~g6065));
assign g22704 = ((~II29372));
assign g30310 = ((~II39773));
assign II17712 = ((~g8031));
assign g27366 = ((~II35686));
assign g17348 = ((~II23436));
assign g11401 = ((~II18359));
assign g25312 = ((~g21211))|((~g14442))|((~g10694))|((~g24590));
assign g19669 = (g1378&g18828);
assign g12055 = ((~g11389));
assign g30610 = ((~g6119)&(~g30412)&(~g25411));
assign g12989 = (g8254&g10273);
assign g5047 = ((~g1264));
assign g20565 = ((~II27020));
assign g10286 = (g6643&g590);
assign II25492 = ((~g18907));
assign II28111 = ((~g20067));
assign g30025 = ((~g29558)&(~g29958));
assign g22030 = ((~g21298)&(~g19557));
assign g24462 = ((~g23803))|((~g3774));
assign g30319 = ((~II39800));
assign g12408 = ((~g11020));
assign II30511 = ((~g21970));
assign g30969 = ((~g30955));
assign g24297 = ((~II31565));
assign g25953 = (g24783&g13699);
assign g21372 = (g9216&g20371);
assign g25252 = ((~g24825)&(~g23680));
assign g5916 = ((~g2309));
assign g29780 = ((~g29480)&(~g29232));
assign II28191 = ((~g19444))|((~II28189));
assign g16817 = ((~II22789));
assign g23423 = (g21602&g22443);
assign II34788 = ((~g26471));
assign g19027 = ((~II25144));
assign g22057 = ((~g21322)&(~g19589));
assign g19677 = (g4182&g17476);
assign II26388 = ((~g17094));
assign II34056 = ((~g25206));
assign g15855 = ((~g13354))|((~g12392));
assign g22025 = ((~g21284)&(~g19549));
assign II40868 = ((~g30740));
assign II24711 = ((~g15296))|((~II24709));
assign g19673 = (g2013&g18829);
assign g21813 = (g20146)|(g20118)|(g18597)|(g19104);
assign g26172 = ((~II34068));
assign g21071 = ((~g19925)&(~g18222));
assign II38355 = ((~g29039));
assign g4803 = ((~g1421));
assign g24107 = ((~g22431));
assign g19328 = (g17098&g8594);
assign g18153 = (g5221&g15704);
assign g26563 = ((~g25530));
assign g11620 = ((~g10601));
assign g27765 = ((~g27552)&(~g27103));
assign g8324 = ((~II15526));
assign g28484 = (g18436&g28177);
assign g9872 = (g6838&g4085);
assign g27278 = ((~g27006)&(~g26319));
assign g21920 = (g5773&g20531);
assign g19670 = (g4156&g17465);
assign II14580 = ((~g2429));
assign g17160 = ((~II23199))|((~II23200));
assign II19479 = ((~g10549));
assign g8045 = ((~g3207));
assign II38609 = ((~g28874));
assign II29972 = ((~g22669));
assign g29414 = ((~II38623));
assign g9203 = ((~g5899));
assign g11833 = ((~g9665)&(~g9780)&(~g9908));
assign g28700 = ((~II37647));
assign g22437 = ((~II28981));
assign g18869 = ((~II24894));
assign g20935 = ((~g19715)&(~g17618));
assign g19534 = ((~g16954));
assign g22720 = ((~g20866))|((~g20956));
assign g15390 = ((~g12279));
assign g3772 = ((~II13224));
assign II30167 = ((~g22598));
assign g18047 = (g5101&g15635);
assign g24537 = ((~g15580)&(~g23899));
assign g24082 = ((~g22887))|((~g14316));
assign g22665 = (g20920&g6153);
assign II29110 = ((~g20738));
assign g24100 = ((~g20885))|((~g22175));
assign g25746 = ((~II33577));
assign g23269 = ((~II30260));
assign g11014 = ((~II17925));
assign g9093 = (g3306&g7676);
assign g10516 = (g7015&g5075);
assign g27051 = ((~g4456)&(~g26081));
assign g30805 = ((~II40667));
assign g23206 = ((~II30071));
assign g17990 = (g5038&g15599);
assign II17813 = ((~g5707));
assign g14467 = ((~g12154));
assign g11558 = ((~II18650));
assign II39411 = ((~g29659));
assign g4029 = ((~g838));
assign g24731 = ((~g23909)&(~g22793));
assign g18484 = ((~II24521))|((~II24522));
assign g25643 = ((~II33466));
assign g25341 = ((~g24923));
assign g30124 = ((~II39635));
assign II30035 = ((~g22705));
assign II26972 = ((~g16913));
assign g20353 = ((~g13702)&(~g16864));
assign g3834 = ((~II13236));
assign g21927 = ((~g20045));
assign g29035 = ((~II37994));
assign g29507 = ((~II38851));
assign g20161 = (g18337&g9426);
assign II18479 = ((~g8820));
assign II16936 = ((~g6100));
assign g21331 = ((~g20472)&(~g16153));
assign g30370 = ((~II39919));
assign g9122 = (g7265&g7763);
assign g5601 = ((~g3092));
assign g5548 = ((~g105));
assign II17843 = ((~g8031));
assign g23769 = (g18048&g23020);
assign II37484 = ((~g27764));
assign II13137 = ((~g33));
assign II34653 = ((~g26165));
assign g23511 = ((~g10714))|((~g14529))|((~g22341));
assign II30275 = ((~g22156));
assign g30782 = ((~II40614));
assign g28118 = ((~II36780))|((~II36781));
assign II22019 = ((~g11731));
assign g4012 = ((~g179));
assign g30860 = ((~II40832));
assign g21851 = ((~g19252)&(~g8842));
assign II23190 = ((~g9507))|((~g13999));
assign g19205 = (g18556)|(g17942);
assign g24595 = (g23502&g23489);
assign g17327 = ((~II23415));
assign g30936 = ((~g30763)&(~g30764));
assign g5948 = ((~g2324));
assign g16633 = ((~II22676));
assign g15188 = ((~g11833));
assign g18542 = ((~II24612))|((~II24613));
assign g13476 = ((~g12565))|((~g3254));
assign g30822 = ((~II40718));
assign g23895 = ((~II31159));
assign g27869 = ((~g27632)&(~g25437));
assign II18326 = ((~g6713));
assign g18873 = ((~g15404));
assign g24133 = ((~g22490));
assign II32925 = ((~g24587));
assign g11854 = ((~g11078));
assign g28047 = ((~II36598));
assign g8168 = ((~g2556));
assign g13613 = ((~II20839));
assign g13374 = ((~g8183)&(~g8045)&(~g11190)&(~g11069));
assign g13895 = ((~g12755));
assign g9232 = ((~g5752));
assign g27218 = ((~II35491));
assign g10309 = (g6783&g4677);
assign g27058 = (g22108&g26624);
assign g9084 = ((~g5848));
assign g16989 = (g6974&g15262);
assign g29527 = (g28748&g29368);
assign g17696 = (g4552&g15360);
assign g24861 = (g24126&g20448);
assign II23398 = ((~g15820));
assign g6301 = ((~g2072));
assign g5996 = ((~g2261));
assign g29061 = ((~II38018));
assign g10831 = ((~g5769)&(~g5817)&(~g5863));
assign g6197 = ((~g3099));
assign g11389 = ((~II18347));
assign g26598 = ((~g25634));
assign II27385 = ((~g19369));
assign II16897 = ((~g6643));
assign g20038 = (g18522&g18464&II26472);
assign II25616 = ((~g1426))|((~g18379));
assign g30617 = ((~g23850)&(~g30412));
assign g23104 = (g20842&g15859);
assign g7328 = ((~g2618));
assign g29702 = ((~II39160));
assign g8302 = ((~II15511));
assign II38728 = ((~g29334));
assign g17648 = ((~g16384));
assign g17235 = ((~g16030)&(~g16047));
assign g16097 = ((~g12837));
assign g7424 = ((~g2633));
assign g19568 = (g8141&g17285);
assign g17390 = ((~II23478));
assign II26240 = (g18174&g18341&g17974);
assign g9319 = (g6369&g8001);
assign g26103 = ((~g25565)&(~g25626));
assign II34444 = ((~g25272));
assign II24657 = ((~g14592))|((~II24655));
assign g12601 = ((~II19747));
assign g8246 = ((~g2978));
assign g29731 = ((~g29583)&(~g1913));
assign II27152 = ((~g20360));
assign g24986 = ((~g23513))|((~g762));
assign II30792 = ((~g14079))|((~II30790));
assign g29085 = ((~II38056));
assign g11962 = ((~g10085)&(~g10173)&(~g10260));
assign II22587 = ((~g14684));
assign g22811 = (g562)|(g559)|(g12451)|(g21851);
assign II38111 = ((~g28371));
assign II23542 = ((~g15835));
assign g22167 = ((~g21446)&(~g19780));
assign g22718 = ((~II29408));
assign g5333 = ((~g2000));
assign g9926 = (g6783&g4168);
assign II21780 = ((~g13305));
assign g22404 = ((~g21631));
assign g25874 = ((~g25085)&(~g21703));
assign II36227 = ((~g27594));
assign g10017 = ((~II16987));
assign g24541 = (g23420&g17896&g23052);
assign II24465 = ((~g14360))|((~II24464));
assign g13268 = ((~g10109));
assign g10416 = ((~II17370));
assign g4188 = ((~g2230));
assign g13836 = ((~g13356));
assign II21395 = ((~g13034));
assign g7052 = ((~II14888));
assign g28657 = (g27925&g13700);
assign g28254 = ((~II37011));
assign g11892 = ((~g11135));
assign g8245 = ((~g2560));
assign g22550 = ((~II29104));
assign g5421 = ((~II13977));
assign g19893 = ((~II26337));
assign II40880 = ((~g30818));
assign g23664 = (g4246&g22552);
assign g19019 = ((~II25120));
assign g12030 = ((~II19211));
assign g17230 = ((~II23314));
assign g29779 = ((~g13943)&(~g29502));
assign g25691 = ((~II33517));
assign g16495 = ((~II22587));
assign g22646 = (g1346&g21514);
assign g18497 = ((~II24545))|((~II24546));
assign g13852 = ((~g13391));
assign II19595 = ((~g10810));
assign g27229 = ((~II35524));
assign II18414 = ((~g6783));
assign g16823 = ((~g5362)&(~g13469));
assign g12828 = ((~g8407)&(~g8447)&(~g8472));
assign g24123 = ((~g22461));
assign g14702 = ((~g11907));
assign g17610 = ((~II23698));
assign II38764 = ((~g29237));
assign g10146 = (g6980&g4386);
assign II36684 = ((~g27317));
assign g29617 = ((~g13989)&(~g29260));
assign g29335 = ((~II38518));
assign g25467 = ((~II33293));
assign II13146 = ((~g42));
assign g26824 = ((~g15491)&(~g26382));
assign II18800 = ((~g11410))|((~II18799));
assign g27359 = (g753&g27010);
assign g13066 = ((~g10872));
assign g20405 = ((~g17585));
assign g4595 = ((~g373));
assign II14634 = ((~g2536));
assign g9480 = (g6574&g8153);
assign II27372 = ((~g19457));
assign g20426 = ((~g17667));
assign g3966 = ((~g1526));
assign II16879 = ((~g4203))|((~g3998));
assign g23580 = ((~II30660));
assign g27950 = ((~g16367)&(~g27673));
assign g13739 = (g7815&g12546);
assign g22632 = (g13992&g21491);
assign g16348 = (g5901&g11983);
assign g6444 = ((~g3102));
assign II14513 = ((~g2190));
assign II29516 = ((~g21020));
assign II30323 = ((~g22799));
assign g19477 = (g14910)|(g16708);
assign g15350 = (g4691&g13201);
assign g19875 = (g14580&g13978&II26317);
assign g26246 = ((~II34192));
assign g27919 = ((~II36382));
assign g22464 = ((~II29010));
assign II24738 = (g14863&g14991&g16266);
assign g5004 = ((~g2516));
assign g22365 = ((~g21192))|((~g21258))|((~g21176));
assign II23633 = ((~g13536));
assign II18088 = ((~g5778));
assign g5797 = (g2406&g2426);
assign g19698 = (g646&g18839);
assign g29089 = ((~II38064));
assign g28719 = (g28482&g19412);
assign g26602 = ((~g25652));
assign g10474 = (g7303&g2661);
assign g18514 = ((~II24566))|((~II24567));
assign g24878 = (g19830&g24210);
assign g7162 = ((~II14920));
assign II33368 = ((~g24444));
assign g30018 = ((~g29533)&(~g29951));
assign g20184 = (g16266&g13764&g13797&II26621);
assign g24545 = ((~g15623)&(~g23910));
assign g23096 = ((~g21178)&(~g19351)&(~g19381));
assign II40002 = ((~g30249));
assign II23782 = ((~g15949));
assign g4061 = ((~g1536));
assign II29663 = ((~g21072));
assign II17792 = ((~g7459));
assign g27882 = ((~g27632)&(~g1220));
assign II40700 = ((~g30648));
assign g22850 = ((~g21858))|((~g21855))|((~g21881));
assign g26488 = (g5301&g25856);
assign II38629 = ((~g29304));
assign II22982 = ((~g15274))|((~II22981));
assign g24851 = ((~II32487));
assign II20410 = ((~g10887));
assign II23104 = ((~g9342))|((~II23103));
assign g12971 = ((~g8526)&(~g8541)&(~g8554));
assign g8823 = ((~II16041));
assign II15244 = ((~g2941))|((~g2944));
assign II40581 = ((~g30703));
assign g30976 = ((~II41102));
assign g30290 = ((~g16459)&(~g29986));
assign g29532 = (g27746&g29372);
assign g18665 = (g14776&g14837&g16189&g13706);
assign II19808 = ((~g8726));
assign g22239 = ((~g20649));
assign II16966 = ((~g4734))|((~II16965));
assign g15547 = ((~II21803));
assign g5358 = ((~g2118));
assign g5855 = ((~g258));
assign g11773 = ((~g9400)&(~g9479)&(~g9603));
assign g24840 = (g9941&g24176);
assign g27001 = (g23364&g26570);
assign II40248 = ((~g30382));
assign g10871 = ((~II17730));
assign g28553 = ((~II37484));
assign g27712 = ((~II36147));
assign g26890 = ((~II35087));
assign g10467 = (g3774&g4994);
assign II40027 = ((~g30253));
assign II14842 = ((~g2214));
assign g12274 = (g7900&g8832);
assign II38770 = ((~g29309));
assign g19885 = (g2746&g18939);
assign II32129 = ((~g24213));
assign g16058 = ((~g6426)&(~g12482)&(~g10952));
assign g8578 = ((~II15784));
assign g22298 = ((~g20760));
assign II30347 = ((~g22872));
assign II35509 = ((~g26836));
assign g26292 = (g4603&g25533);
assign g15777 = ((~II22025));
assign g17297 = ((~II23383));
assign g9603 = (g3566&g8224);
assign g18937 = ((~II24973));
assign II28541 = ((~g21467));
assign g26021 = ((~II33915));
assign g26685 = ((~II34662));
assign g22037 = ((~g21304)&(~g19564));
assign g23364 = ((~g21987))|((~g21981));
assign II14981 = ((~g2625));
assign g27928 = ((~II36393));
assign g30834 = ((~II40754));
assign II37924 = ((~g28529));
assign II32510 = ((~g17815))|((~II32509));
assign II22515 = ((~g13620));
assign II31514 = ((~g23614));
assign g26164 = ((~II34056));
assign II35837 = ((~g26911));
assign g11564 = ((~II18668));
assign g23071 = (g21808)|(g21802)|(g21846);
assign II18338 = ((~g6574));
assign g18643 = ((~g16337));
assign g15052 = ((~II21407));
assign g10851 = ((~g5828)&(~g5873)&(~g5910));
assign g24051 = ((~II31266));
assign II36129 = ((~g27542));
assign g13657 = ((~g12452));
assign g25105 = ((~g23839));
assign g14454 = ((~g12991));
assign g28924 = ((~II37891));
assign II25486 = ((~g18754));
assign II21878 = ((~g11719));
assign g11471 = ((~II18435));
assign II38843 = ((~g15981))|((~II38841));
assign II27047 = ((~g19258));
assign g23838 = ((~II31074));
assign g27509 = (g23945&g27148);
assign g16388 = (g5935&g12039);
assign g12439 = ((~II19595));
assign g22315 = ((~g20786));
assign II32527 = ((~g18038))|((~II32526));
assign II27288 = ((~g19457));
assign g30031 = ((~g24695)&(~g29925));
assign g15271 = ((~II21554));
assign g28369 = ((~II37266));
assign II31610 = ((~g23576));
assign II34327 = ((~g25260));
assign g27261 = ((~g26980)&(~g26263));
assign g9636 = (II16735&II16736);
assign g25612 = ((~II33437));
assign g24410 = ((~II31904));
assign g27686 = ((~II36069));
assign II24103 = ((~g6363))|((~II24102));
assign g24350 = ((~II31724));
assign g25318 = (g24682&g19358&g19335);
assign g20574 = ((~II27047));
assign g28662 = (g27911&g11951);
assign g11546 = ((~II18614));
assign g27801 = ((~II36257))|((~II36258));
assign g29419 = ((~II38638));
assign II28467 = ((~g20942));
assign g8144 = ((~g836));
assign g16467 = ((~II22503));
assign g27282 = ((~g27016)&(~g26332));
assign II38638 = ((~g29311));
assign g8516 = (g6314&g198);
assign g29718 = ((~g6104)&(~g29583)&(~g25409));
assign g19572 = (g8161&g17297);
assign g22170 = ((~g21453)&(~g19788));
assign g21134 = ((~g20111)&(~g20134)&(~g20157));
assign g5009 = ((~g2781));
assign g24564 = (g23435&g18124&g23084);
assign g16832 = ((~II22803));
assign II14472 = ((~g3080));
assign g9961 = ((~g5615));
assign g25771 = ((~g24607));
assign g8972 = (g3650&g1877);
assign g5319 = ((~g2688));
assign g9940 = (g7230&g4179);
assign g11111 = ((~II18025));
assign II20520 = ((~g13246));
assign g26720 = ((~II34767));
assign g28409 = ((~g24676)&(~g27801));
assign g23184 = ((~II30005));
assign II33846 = ((~g25780));
assign g3972 = ((~g1533));
assign II35983 = ((~g26827));
assign II27086 = ((~g19229));
assign g19325 = ((~II25701))|((~II25702));
assign g19519 = ((~g16794));
assign g28833 = ((~II37796));
assign II25866 = ((~g2142))|((~II25865));
assign II18191 = ((~g7922))|((~II18190));
assign g12867 = ((~g8912));
assign g29429 = ((~II38668));
assign g8507 = (g6369&g954);
assign g28037 = ((~II36568));
assign g18355 = ((~II24368));
assign II37653 = ((~g28359));
assign g9354 = ((~II16569));
assign g9245 = ((~II16507));
assign g10929 = ((~g5952));
assign II37080 = ((~g28085));
assign g5967 = ((~g1567));
assign g22788 = (g14454&g21640);
assign g22226 = ((~II28792));
assign g30111 = (g29869&g11425);
assign g21199 = ((~II27766));
assign II32688 = ((~g24028))|((~II32686));
assign g6135 = ((~II14650));
assign g20666 = ((~II27257));
assign II36879 = ((~g27972));
assign II20050 = ((~g10095))|((~II20048));
assign g13970 = (g7655&g12892);
assign g14956 = (g11059&g13151);
assign g8580 = ((~g6281));
assign g13291 = (g5656&g11154);
assign II35072 = ((~g26661));
assign g30796 = ((~g16069)&(~g30696));
assign II19727 = ((~g8726));
assign g30483 = ((~II40059));
assign II30589 = ((~g23133));
assign g22339 = ((~g14442))|((~g21149))|((~g10694));
assign g4156 = ((~g1532));
assign II38042 = ((~g28584));
assign g17813 = (g4757&g15464);
assign g7556 = ((~g1183));
assign g9622 = (g6838&g8239);
assign g11144 = ((~II18058));
assign g26541 = ((~g13755)&(~g25269));
assign II28742 = ((~g21890))|((~II28741));
assign g13643 = (g5431&g12502);
assign g9035 = ((~II16354));
assign g25262 = ((~g24869)&(~g17824));
assign g11521 = ((~II18539));
assign II32538 = ((~g18247))|((~g24080));
assign II19637 = ((~g10872));
assign II17641 = ((~g6215));
assign g11817 = ((~g11008));
assign g7606 = ((~g2190));
assign g21931 = (g4632&g20539);
assign g6427 = ((~g2026));
assign g13459 = ((~II20676));
assign II34921 = ((~g26217));
assign g23029 = ((~g21111)&(~g19267));
assign g24494 = ((~g23716)&(~g23763));
assign g16199 = (g5763&g11867);
assign g10694 = ((~g4326));
assign II29490 = ((~g21009));
assign g12151 = ((~g10374)&(~g10440)&(~g10498));
assign II30496 = ((~g23137));
assign g24839 = ((~II32452))|((~II32453));
assign g15171 = (g8015&g12647);
assign g24395 = ((~II31859));
assign g9902 = (g6912&g4118);
assign II28013 = ((~g19987));
assign g10482 = ((~II17433));
assign g14395 = ((~g12107));
assign g27450 = ((~g26902)&(~g24613));
assign g21486 = (g6832&g20449);
assign g27070 = (g22009&g26631);
assign g15581 = (g5122&g13243);
assign g29929 = ((~g29673)&(~g22367));
assign g14113 = (g7715&g12950);
assign II25821 = ((~g18509))|((~II25819));
assign II26220 = ((~g17691));
assign g6896 = ((~g2824));
assign II16984 = ((~g7936));
assign g29649 = ((~II39065));
assign g26099 = ((~g6068)&(~g24183)&(~g25313));
assign II29432 = ((~g20991));
assign II32324 = ((~g17927))|((~II32323));
assign g28397 = ((~g27869)&(~g22344));
assign g24929 = ((~g23511));
assign g13672 = (g7788&g12522);
assign g7757 = ((~g1701));
assign II25539 = ((~g92))|((~g18174));
assign g23060 = ((~g21606));
assign g18447 = ((~g16120)&(~g14371));
assign II33418 = ((~g25022));
assign g8469 = ((~II15671));
assign II31532 = ((~g23685));
assign g26868 = ((~II35049));
assign g11790 = ((~g9497)&(~g9621)&(~g9745));
assign g26729 = ((~II34794));
assign g24912 = ((~g23495));
assign II31925 = ((~g23469));
assign g26339 = (g4780&g25599);
assign g24206 = ((~g16966)&(~g22228));
assign g22344 = ((~g21233));
assign g12178 = ((~g8378));
assign g30446 = ((~II40002));
assign g11806 = ((~g9582)&(~g9661)&(~g9776));
assign II18838 = ((~g10871));
assign II30242 = ((~g22867));
assign g10311 = (g7015&g4685);
assign g30303 = ((~g13516)&(~g30005));
assign g15721 = ((~g12565))|((~g6314));
assign g23521 = ((~g22920))|((~g14618))|((~g10754));
assign g29030 = ((~g9203))|((~g28540));
assign g8863 = ((~II16117));
assign g24361 = ((~II31757));
assign II40504 = ((~g30683));
assign g29212 = ((~g15219)&(~g28944));
assign g10133 = (g3554&g7162);
assign II18253 = ((~g6783));
assign II25865 = ((~g2142))|((~g18573));
assign II31235 = ((~g22218));
assign g26046 = ((~g25618)&(~g24899));
assign g9465 = ((~II16641));
assign II37778 = ((~g28567));
assign g10660 = (g3650&g1991);
assign II34974 = ((~g26168));
assign g27206 = ((~II35455));
assign g26804 = ((~g15172)&(~g26235));
assign g4898 = ((~g605));
assign g21966 = ((~II28524));
assign g12642 = ((~g8771));
assign g8940 = ((~II16238));
assign g7149 = ((~g3105));
assign g13461 = ((~II20682));
assign g27155 = ((~g26434));
assign g16999 = (g7224&g15354);
assign II35011 = ((~g26304));
assign II37089 = ((~g28103));
assign g19622 = ((~II26051));
assign g17129 = (g8079&g15679);
assign g28343 = ((~II37232));
assign g22087 = ((~g21349)&(~g19630));
assign g13588 = ((~II20810));
assign g16854 = ((~g15802)&(~g13010));
assign g23502 = ((~g22879))|((~g14529))|((~g10714));
assign g25115 = ((~g23879));
assign g30330 = (g30195&g8333);
assign g20918 = ((~g19687)&(~g17554));
assign II25596 = ((~g61))|((~II25595));
assign g30492 = (g30187&g11414);
assign g13137 = ((~g9822))|((~g7358));
assign II40697 = ((~g30647));
assign g8239 = ((~g2221));
assign g16990 = (g7912&g15306);
assign g9629 = ((~II16726));
assign g23486 = ((~g22844))|((~g14442))|((~g10694));
assign g25322 = ((~g24883));
assign II15827 = ((~g3806));
assign g21576 = (g19067)|(g16924)|(g14301);
assign g15719 = ((~g13401))|((~g12392));
assign g21233 = ((~g19418)&(~g17145));
assign g30815 = ((~II40697));
assign g26449 = (g5201&g25802);
assign g27660 = (g26835&g11117);
assign g25862 = ((~II33708));
assign II36490 = ((~g27265));
assign II41041 = ((~g30801));
assign g8164 = ((~g2562));
assign II33567 = ((~g25049));
assign II29148 = ((~g20892));
assign II15451 = ((~g3238));
assign II24704 = ((~g14554))|((~II24702));
assign g13313 = ((~g8183)&(~g11332)&(~g11190)&(~g7880));
assign g18822 = ((~g15179));
assign g29174 = (g29031&g20684);
assign g11732 = ((~g10826));
assign g12185 = ((~g10415)&(~g10478)&(~g10539));
assign g5289 = ((~g2808));
assign II38686 = ((~g29316));
assign g22840 = ((~II29641));
assign g29822 = (g29705&g22335);
assign g17363 = ((~II23451));
assign g19545 = (g16943&g16791&g14863);
assign g30827 = ((~II40733));
assign g23440 = (g22870&g19680);
assign g5610 = ((~g1476));
assign g26036 = (g25413&g19502);
assign II17762 = ((~g7333));
assign g23527 = (g5905&g22353);
assign g9610 = ((~II16714));
assign g27106 = ((~g4985)&(~g26103));
assign g17868 = ((~II23929));
assign g12377 = (g7553)|(g11059);
assign g28608 = ((~g27831));
assign g10037 = (g6678&g4231);
assign g11952 = ((~g10065)&(~g10156)&(~g10226));
assign II15925 = ((~g6751));
assign g27532 = ((~g26761)&(~g25182));
assign g11617 = ((~g8313))|((~g2883));
assign II30832 = ((~g22099));
assign g12049 = ((~g10220)&(~g10306)&(~g10384));
assign II36554 = ((~g27283));
assign g20535 = ((~g18523));
assign g28030 = ((~II36551));
assign g11154 = ((~II18070));
assign II20661 = ((~g12442));
assign g23537 = ((~g10754))|((~g14618))|((~g22384));
assign g4778 = ((~g1131));
assign II38665 = ((~g29412));
assign g26780 = (g26119&g16622);
assign g5372 = ((~g2119));
assign g19915 = ((~II26365));
assign II25665 = ((~g2120))|((~II25664));
assign g23296 = ((~II30341));
assign g21052 = ((~g19900)&(~g18106));
assign g28028 = (g27595&g9898);
assign g3963 = ((~g863));
assign g30437 = (g30139&g11082);
assign g11851 = (g7849&g8670);
assign g16067 = (g7700&g11774);
assign g26827 = ((~g15577)&(~g26425));
assign II21641 = ((~g13068));
assign g26092 = ((~II33990));
assign g11585 = ((~II18731));
assign g30345 = (g30195&g8388);
assign II17740 = ((~g8031));
assign g21658 = (g2896&g20501);
assign II23409 = ((~g15822));
assign g17598 = (g4380&g15265);
assign g8437 = (g3410&g915);
assign g16139 = (g5704&g11824);
assign g16073 = (g5605&g11778);
assign g5974 = ((~g2327));
assign g29150 = ((~II38193));
assign g26833 = (g5651&g26237);
assign II37813 = ((~g28388))|((~g28391));
assign g18333 = (g2888&g15777);
assign g24956 = ((~II32716));
assign g8025 = ((~g3050));
assign g6363 = ((~g653));
assign II15487 = ((~g3250));
assign g15872 = ((~g12711))|((~g7085));
assign g22076 = ((~g21340)&(~g19619));
assign g29443 = ((~II38710));
assign II27303 = ((~g19369));
assign II38097 = ((~g28364));
assign g23444 = ((~g22945));
assign g29962 = (g29789&g29069);
assign g24795 = (g12017&g24232);
assign II28076 = ((~g20025));
assign II29402 = ((~g20978));
assign II40518 = ((~g30688));
assign g19601 = (g640&g18784);
assign g6035 = ((~g2165));
assign g18785 = ((~g15040));
assign g7595 = ((~g2900));
assign g26131 = ((~II34026));
assign g17838 = (g4803&g15488);
assign g30257 = ((~g16290)&(~g30091));
assign II16354 = ((~g3618));
assign II35059 = ((~g26126))|((~II35057));
assign g20881 = ((~g19603)&(~g17398));
assign g23142 = ((~g21825));
assign II29993 = ((~g22704));
assign II28833 = ((~g21470));
assign g15707 = ((~II21955));
assign g19102 = (g15003&g18796&g16325&g16371);
assign g13561 = ((~g12657))|((~g3566));
assign g30395 = (g30241&g9000);
assign g26805 = ((~g15173)&(~g26236));
assign g19715 = (g2013&g18845);
assign II36483 = ((~g27264));
assign g14144 = ((~II21096));
assign g7796 = ((~g1008));
assign g11574 = ((~II18698));
assign II40844 = ((~g30823));
assign g12171 = ((~g10398)&(~g10461)&(~g10522));
assign g5943 = ((~g1918));
assign g17220 = ((~g15962)&(~g14703));
assign g15901 = ((~g12711))|((~g7085));
assign g8534 = (g3410&g879);
assign g12308 = ((~g8312));
assign g21877 = ((~g18611))|((~g19246))|((~g19257));
assign g26361 = (g4888&g25637);
assign g16219 = (g8295&g11878);
assign g30360 = ((~II39895));
assign II35057 = ((~g26137))|((~g26126));
assign II19530 = ((~g10653));
assign g27847 = ((~II36321));
assign g10793 = ((~g5658)&(~g5687)&(~g5728));
assign g21945 = ((~II28461));
assign g17600 = (g4386&g15271);
assign g16163 = (g5736&g11841);
assign g6156 = ((~II14668));
assign g6141 = ((~g554));
assign II19380 = ((~g10606));
assign II38077 = ((~g28357));
assign II26714 = ((~g17720));
assign g30947 = (g30936&g20760);
assign g18388 = ((~g14486));
assign II33466 = ((~g25053));
assign g12331 = (g7927&g8882);
assign II18767 = ((~g10086));
assign g30571 = ((~g30401));
assign II30816 = ((~g22092));
assign g17176 = (g7742&g14298);
assign g19561 = (g8068&g17262);
assign g11698 = ((~g9676))|((~g3522));
assign II34183 = ((~g25241));
assign g26676 = ((~g25377)&(~g17181));
assign g27211 = ((~II35470));
assign g27285 = ((~g27019)&(~g26339));
assign g7615 = ((~g3123));
assign g25811 = ((~II33649));
assign g5709 = (g337&g368);
assign g22195 = ((~g21527)&(~g19859));
assign g7592 = ((~g2540));
assign g21015 = ((~g19846)&(~g17924));
assign g23634 = ((~II30766));
assign g22443 = ((~g21036));
assign g10273 = ((~II17235));
assign II16079 = ((~g6086));
assign g4047 = ((~g1095));
assign g30881 = ((~II40895));
assign II30686 = ((~g23136));
assign g29258 = ((~II38369));
assign g12598 = ((~g8757));
assign g11456 = ((~II18420));
assign II32901 = ((~g25121));
assign II40823 = ((~g30806));
assign g29233 = (g9374&g28799);
assign g20272 = (g18708&g18789&g13724&g16395);
assign g28236 = ((~II36957));
assign g29210 = ((~g28919)&(~g28462));
assign g29287 = ((~g28810));
assign g22772 = ((~II29530));
assign g19860 = (g2720&g18923);
assign g30848 = ((~II40796));
assign g5863 = (g1024&g1011);
assign g7971 = ((~g3049));
assign g6678 = ((~II14811));
assign g28388 = ((~II37312))|((~II37313));
assign g14472 = ((~g12992));
assign g15763 = ((~g12657))|((~g6783));
assign g19608 = ((~g16913));
assign g28495 = ((~g27244)&(~g27723));
assign g26914 = ((~g26107)&(~g22319));
assign g25661 = ((~II33485));
assign II41120 = ((~g30978));
assign g21305 = (g9232&g20297);
assign g12967 = ((~g8517)&(~g8532)&(~g8546));
assign g17962 = ((~II23999));
assign g8905 = ((~II16185));
assign g8630 = ((~II15818));
assign g29640 = ((~II39038));
assign g28951 = ((~II37920));
assign II21482 = ((~g13058));
assign II25246 = ((~g17233));
assign g22230 = ((~g20634));
assign II30116 = ((~g22762));
assign g29942 = (g29771&g28877);
assign g25626 = (g24504&g17865);
assign g23578 = (g3960&g22458);
assign II28443 = ((~g19358));
assign g11821 = ((~g10848));
assign g28302 = ((~II37155));
assign g22255 = (g21661&g12242);
assign g20672 = ((~g20164))|((~g3254));
assign g10383 = (g6980&g4794);
assign II30707 = ((~g22059));
assign g22670 = ((~II29304));
assign g23739 = ((~II30931));
assign g28723 = ((~g28528));
assign g16743 = ((~g14936));
assign g18885 = ((~g13847)&(~g12129));
assign II32647 = ((~g24093))|((~II32645));
assign g6572 = ((~g972));
assign g15228 = ((~II21511));
assign g9009 = (g6486&g565);
assign g30778 = ((~II40600));
assign g8277 = ((~g3305));
assign g27436 = ((~g23118)&(~g27187)&(~g24427));
assign g17158 = ((~II23191))|((~II23192));
assign g30757 = (g30601&g20780);
assign g25976 = ((~II33790));
assign g13021 = ((~g9534))|((~g6912));
assign II32388 = ((~g23385));
assign II18121 = ((~g3254));
assign g29804 = ((~II39264));
assign g24599 = ((~II32181));
assign II23539 = ((~g13524));
assign g24150 = ((~g22527));
assign g24616 = ((~g499))|((~g23376));
assign g11939 = ((~g10041)&(~g10116)&(~g10206));
assign II29635 = ((~g21062));
assign g15287 = ((~II21563));
assign II18389 = ((~g6519));
assign g25993 = ((~II33831));
assign g19143 = (g17174&g16761);
assign g25164 = ((~II32970));
assign g22201 = (g21271&g16881);
assign g18464 = ((~II24494))|((~II24495));
assign II22901 = ((~g15022))|((~II22900));
assign g30246 = ((~g16107)&(~g30079));
assign g24275 = ((~II31499));
assign g20375 = ((~g13739)&(~g16879));
assign g23282 = ((~II30299));
assign II17721 = ((~g6641));
assign II16363 = ((~g3900));
assign g23940 = ((~g22376));
assign g29566 = (g26047&g29395);
assign g23616 = (g17724&g22988);
assign g16447 = (g5983&g12147);
assign II31027 = ((~g22155));
assign g10528 = (g7265&g5107);
assign g13869 = ((~g11638));
assign II18268 = ((~g7085));
assign g8925 = ((~II16215));
assign g10197 = (g6448&g441);
assign II33476 = ((~g24453));
assign II41017 = ((~g30768))|((~g30771));
assign II31062 = ((~g23003));
assign II25977 = ((~g16692));
assign g8845 = ((~II16085));
assign II37702 = ((~g28512));
assign g17123 = ((~II23132))|((~II23133));
assign g20370 = ((~g17468));
assign g21907 = ((~g19972));
assign g22624 = (g13983&g21483);
assign g20000 = (g18449&g18369&II26440);
assign g6117 = ((~II14634));
assign II16312 = ((~g5424));
assign g30987 = ((~II41135));
assign g17984 = ((~g14008));
assign II41010 = ((~g30775))|((~g30779));
assign g16381 = (g5926&g12021);
assign g16622 = ((~II22667));
assign g20945 = ((~g19732)&(~g17653));
assign g13483 = (g6020&g12209);
assign II23045 = ((~g9248))|((~g13894));
assign g17902 = (g4905&g15534);
assign g27132 = ((~II35319));
assign g19413 = (g16954&g16602&g14507);
assign II18671 = ((~g8812));
assign g7733 = ((~g1007));
assign g27192 = ((~II35413));
assign g25197 = ((~g24528)&(~g10340));
assign g25452 = ((~g16101)&(~g25117));
assign g13506 = (g5921&g11638);
assign g25061 = ((~g23803))|((~g7265));
assign II31712 = ((~g23890));
assign g21111 = (g19524&g14395&g16529);
assign II27253 = ((~g19420));
assign g28478 = (g18358&g28175);
assign g27554 = (g24004&g27164);
assign g19305 = ((~g16626));
assign g5821 = ((~g1600));
assign g21177 = (g5865&g19309);
assign g13367 = ((~II20458));
assign g20591 = ((~II27098));
assign g19400 = ((~II25820))|((~II25821));
assign g21900 = (g19306&g13011);
assign II28953 = ((~g21659));
assign g17966 = (g5012&g15585);
assign g13270 = (g985&g11102);
assign g26696 = ((~II34695));
assign II28500 = ((~g21457));
assign g17487 = ((~II23575));
assign II32498 = ((~g18155))|((~g24069));
assign g23916 = ((~II31188));
assign II23857 = ((~g13560));
assign g28200 = ((~II36864));
assign g25668 = ((~g20858)&(~g24437));
assign g5196 = ((~g2114));
assign g6085 = ((~II14602));
assign g12565 = ((~II19739));
assign g12854 = ((~II19915));
assign g22448 = ((~II28994));
assign g27348 = ((~g27109)&(~g26494));
assign II41066 = ((~g30926))|((~II41064));
assign g19790 = (g4564&g17704);
assign g12156 = ((~g8344));
assign II18094 = ((~g7085));
assign g7849 = ((~g2956));
assign g21394 = (g9216&g20390);
assign g9382 = (g6519&g8065);
assign g28191 = ((~g27365)&(~g26860));
assign g24805 = ((~II32365));
assign g21496 = ((~II28034));
assign gbuf107 = (g1260);
assign g20478 = ((~II26923));
assign g30592 = ((~II40320));
assign g5218 = ((~g2787));
assign g29310 = (g28978&g28951);
assign g15941 = ((~g12657))|((~g6574));
assign g6028 = ((~g2345));
assign II35440 = ((~g27186));
assign II16633 = ((~g6486));
assign II29736 = ((~g20884));
assign g27916 = ((~g16219)&(~g27659));
assign g30891 = ((~II40925));
assign g15502 = ((~II21761));
assign g17475 = (g4179&g15148);
assign g29954 = (g29770&g28975);
assign g21192 = (g19419&g19400&II27755);
assign g21980 = ((~g21252)&(~g19531)&(~g19540));
assign g29207 = ((~g28914)&(~g28460));
assign II25532 = ((~g52))|((~g18179));
assign II24625 = ((~g6136))|((~II24624));
assign II31257 = ((~g22234));
assign g5075 = ((~g1769));
assign g25296 = ((~II33128));
assign II37098 = ((~g27918));
assign g18597 = (g13714&g13791&II24689);
assign II32586 = ((~g17815))|((~g23937));
assign g27074 = (g22118&g26635);
assign g7655 = ((~g1002));
assign g6173 = ((~g557));
assign g10126 = ((~II17100));
assign g18846 = ((~g15290));
assign g18573 = ((~g14596));
assign g9531 = ((~II16684));
assign gbuf2 = (g2861);
assign g22251 = ((~g20666));
assign g23076 = ((~g17023)&(~g21129));
assign g30439 = ((~II39991));
assign g18436 = ((~g14454));
assign g10508 = (g6751&g5053);
assign g22050 = ((~g19450))|((~g21244))|((~g19503));
assign II39764 = ((~g30060));
assign gbuf184 = (g2417);
assign g5883 = (g2406&g2456);
assign g12688 = ((~g8794));
assign g22116 = ((~g21374)&(~g19678));
assign g30799 = ((~II40651));
assign g27924 = (g13983&g27422);
assign g27173 = ((~g26490));
assign g30560 = ((~II40260));
assign g28040 = ((~II36577));
assign II39889 = ((~g30285));
assign g26270 = (g25903&g9465);
assign II22569 = ((~g14955));
assign g11970 = ((~g11271));
assign g13849 = ((~g13381));
assign g23614 = ((~II30728));
assign g10779 = ((~II17627));
assign II34901 = ((~g26295));
assign g9049 = (g5473&g7619);
assign g13004 = (g10186&g8317);
assign g30514 = ((~II40122));
assign g27965 = ((~II36432));
assign g10454 = (g3618&g1825);
assign g29662 = ((~g29570));
assign II23602 = ((~g13529));
assign II37305 = ((~g27900))|((~II37303));
assign g24419 = ((~II31931));
assign g27629 = ((~g26829)&(~g26051));
assign g10462 = (g7230&g4970);
assign II18602 = ((~g9591));
assign g11300 = ((~II18250));
assign g23596 = ((~II30692));
assign g10062 = (g3566&g4275);
assign II33377 = ((~g25033));
assign g24847 = ((~g16356)&(~g24247));
assign II20799 = ((~g13155));
assign g28454 = (g26121&g28167);
assign g30256 = ((~g16282)&(~g30090));
assign II25064 = ((~g14395));
assign II18467 = ((~g8769));
assign g29479 = (g21461&g29280);
assign g30271 = ((~g16388)&(~g30105));
assign g27945 = (g4376&g27451);
assign II29660 = ((~g21071));
assign g20954 = ((~g19753)&(~g17696));
assign g13211 = ((~g9730));
assign g10537 = (g7488&g5126);
assign g22677 = ((~II29323));
assign g22042 = ((~g21309)&(~g19569));
assign g18907 = ((~g14336)&(~g12429));
assign II23019 = ((~g9216))|((~II23018));
assign g13926 = ((~g11832));
assign g22415 = ((~II28959));
assign g29077 = ((~II38042));
assign g27576 = ((~II35993))|((~II35994));
assign II29519 = ((~g21021));
assign g27245 = (g26877&g22286);
assign II23967 = ((~g14092))|((~II23966));
assign g20580 = ((~II27065));
assign g27302 = ((~g27042)&(~g26379));
assign II18668 = ((~g8756));
assign II39246 = ((~g29692));
assign II21736 = ((~g11702));
assign II38827 = ((~g29355));
assign g22795 = ((~II29569));
assign II31592 = ((~g23553));
assign II23010 = ((~g13926))|((~II23008));
assign g19481 = ((~g16629));
assign g12949 = ((~g8510)&(~g8525)&(~g8540));
assign g23114 = ((~g17114)&(~g21181));
assign g19775 = (g1346&g18875);
assign g13203 = ((~g9623));
assign g16092 = ((~g12830));
assign g29377 = ((~g28967));
assign g27409 = (g1378&g27137);
assign g20149 = (g13764&g13797&II26599);
assign II17103 = ((~g3494));
assign II20466 = ((~g11330))|((~II20465));
assign g10153 = (g6574&g4398);
assign g7455 = ((~g2740));
assign II16244 = ((~g5416));
assign g7868 = ((~g2584));
assign g28109 = ((~II36758));
assign II40841 = ((~g30817));
assign g26238 = ((~II34180));
assign II35389 = ((~g26168));
assign g13114 = ((~g9676))|((~g6980));
assign g23801 = ((~II31027));
assign g26356 = ((~g16539))|((~g25183));
assign II40871 = ((~g30746));
assign g29359 = ((~II38548));
assign g26265 = ((~g25972)&(~g13360));
assign g10530 = (g3774&g2519);
assign g23546 = ((~II30594));
assign g30252 = ((~g16217)&(~g30086));
assign g29997 = (g29918&g22277);
assign g11670 = ((~II18854));
assign II33307 = ((~g25011));
assign II20278 = ((~g9027));
assign II35449 = ((~g27154));
assign g26212 = (g4217&g25467);
assign g11422 = ((~II18386));
assign g10912 = ((~II17795));
assign II16723 = ((~g5556));
assign II27179 = ((~g20419));
assign II33300 = ((~g25112));
assign g20044 = (g5375&g18539);
assign g23175 = ((~II29978));
assign g15418 = ((~II21680));
assign g19013 = ((~II25102));
assign g19977 = ((~g18630));
assign II22699 = ((~g14677));
assign g28067 = ((~II36644));
assign g11885 = (g7834&g8684);
assign g28384 = ((~II37296))|((~II37297));
assign g19616 = (g3966&g17363);
assign g10582 = (g7053&g5182);
assign g26343 = (g4821&g25609);
assign II34009 = ((~g25882));
assign g7975 = ((~g39));
assign II39840 = ((~g30272));
assign II40066 = ((~g30260));
assign II18539 = ((~g11290));
assign II34731 = ((~g26341));
assign g10908 = ((~II17783));
assign g12930 = ((~g8493)&(~g8509)&(~g8524));
assign g22138 = ((~g21396)&(~g19718));
assign II25315 = ((~g16895));
assign g10557 = (g6643&g617);
assign g4363 = ((~g821));
assign g10376 = (g3494&g1259);
assign g29435 = ((~II38686));
assign g16242 = (g5806&g11893);
assign g13284 = ((~g10179));
assign g29516 = ((~II38878));
assign g15379 = ((~II21641));
assign II30200 = ((~g22740));
assign g20618 = ((~II27179));
assign g21971 = ((~g21243)&(~g19499));
assign g20749 = ((~II27338));
assign g26928 = ((~g25781))|((~g26374))|((~g25725));
assign II23244 = ((~g13882))|((~II23242));
assign II39976 = ((~g30245));
assign g18976 = ((~g15777));
assign II38671 = ((~g29171));
assign g22279 = ((~g20725));
assign g27505 = ((~II35863));
assign g13513 = (g6043&g12289);
assign g25919 = ((~g24973));
assign g28444 = (g28137&g9273);
assign g21043 = ((~g19884)&(~g18058));
assign g4412 = ((~g2083));
assign g5752 = ((~g113));
assign g22827 = ((~II29610));
assign g25707 = ((~II33535));
assign II36117 = ((~g27539));
assign II30293 = ((~g22693));
assign II14584 = ((~g465));
assign g27220 = ((~II35497));
assign g28325 = ((~g27747)&(~g10238));
assign II21514 = ((~g13041));
assign g8096 = ((~II15359));
assign II36966 = ((~g28012));
assign g20158 = (g18543&g9886);
assign g23853 = ((~g22300));
assign g22455 = ((~II29001));
assign g20465 = ((~g17862));
assign g22243 = ((~II28813));
assign g29497 = ((~II38807));
assign gbuf100 = (g1231);
assign g22765 = ((~II29513));
assign g15402 = (g4620&g12783);
assign g21976 = ((~g19242))|((~g21120))|((~g19275));
assign g8977 = ((~II16289));
assign II27197 = ((~g20459));
assign II18656 = ((~g8872));
assign g8882 = ((~II16150));
assign g28004 = ((~II36493));
assign g30545 = ((~II40215));
assign g20191 = (g18543&g9758);
assign g15833 = ((~g12565))|((~g6314));
assign II38916 = ((~g29201));
assign g5696 = (g1706&g1730);
assign g27698 = ((~II36105));
assign g19154 = ((~g17382)&(~g15094));
assign g19090 = (g18744&g15080&g13774&g16371);
assign II31050 = ((~g22162));
assign g16213 = ((~g12249));
assign g9673 = ((~II16766));
assign g26931 = ((~g25861))|((~g26417))|((~g25798))|((~g25835));
assign II22823 = ((~g13613));
assign g26918 = ((~g25826))|((~g26374))|((~g25725))|((~g25781));
assign g19179 = ((~g17719)&(~g15453));
assign g27691 = ((~II36084));
assign g30877 = ((~II40883));
assign g10905 = ((~g5923));
assign II18813 = ((~g10850));
assign g26786 = ((~g26049)&(~g22777));
assign g15849 = ((~g12657))|((~g6783));
assign II37620 = ((~g28611));
assign g30640 = ((~g16187)&(~g30437));
assign g30447 = (g30143&g11145);
assign g20393 = ((~g17548));
assign g22636 = ((~II29238));
assign g20729 = ((~II27318));
assign g27550 = ((~II35945))|((~II35946));
assign g14537 = ((~g12208));
assign g20277 = (g13805&g13825&II26690);
assign II22317 = ((~g2934))|((~II22316));
assign II19318 = ((~g10486));
assign II36766 = ((~g27339));
assign II31880 = ((~g23799));
assign g13090 = ((~g9676))|((~g6980));
assign II35876 = ((~g26813));
assign g12470 = ((~II19654));
assign gbuf205 = (g2648);
assign g19694 = (g4211&g17493);
assign g10593 = (g7303&g5213);
assign II16521 = ((~g5512));
assign g22124 = ((~g21380)&(~g19694));
assign II20658 = ((~g11845));
assign g29461 = ((~II38764));
assign g30535 = ((~II40185));
assign g20912 = ((~g19668)&(~g17529));
assign g12175 = ((~g8369));
assign g7078 = ((~g1924));
assign g17302 = ((~g16103)&(~g16135));
assign g29741 = ((~g6104)&(~g29583)&(~g25376));
assign g21454 = (g9277&g20435);
assign g4246 = ((~g865));
assign g27257 = ((~g26971)&(~g26243));
assign g10747 = ((~g3866))|((~g7488));
assign g27125 = ((~g26451))|((~g7265));
assign II37875 = ((~g28501));
assign g20159 = (g16809&g9288);
assign II21655 = ((~g11696));
assign g14601 = ((~g12268));
assign g22155 = ((~g21425)&(~g19757));
assign g24166 = ((~g22570));
assign II39550 = ((~g29848));
assign g13840 = ((~g12455));
assign g10364 = (g6486&g4749);
assign II19545 = ((~g10617));
assign II39267 = ((~g29702));
assign g23685 = ((~II30847));
assign g9061 = (g3306&g7623);
assign g7679 = ((~g1003));
assign g26836 = ((~II34977));
assign II22707 = ((~g15661))|((~II22705));
assign g29482 = (g21461&g29285);
assign II33198 = ((~g25067));
assign II16144 = ((~g6101));
assign g7347 = ((~g490));
assign g26042 = ((~g25505)&(~g24867));
assign g14849 = ((~g12152));
assign g12045 = ((~II19226));
assign II24227 = ((~g6427))|((~II24226));
assign g18522 = ((~II24576))|((~II24577));
assign II26481 = ((~g18590));
assign g13323 = ((~II20390));
assign II40682 = ((~g30642));
assign g6183 = ((~g291));
assign II32120 = ((~g24209));
assign g24653 = (g24095)|(g20850);
assign g30957 = ((~g30920)&(~g30947));
assign II31871 = ((~g23765));
assign II29405 = ((~g20979));
assign II39472 = ((~g29937));
assign g19031 = ((~II25156));
assign II34192 = ((~g25243));
assign g12544 = ((~g8305))|((~g5556));
assign g29463 = ((~II38770));
assign g18982 = (g13519&g16154);
assign g10858 = ((~II17709));
assign g27700 = ((~II36111));
assign g19547 = (g16943&g16770&g14922);
assign II21119 = ((~g12523));
assign g11332 = ((~g4094));
assign II38369 = ((~g29112));
assign g24232 = ((~g22637)&(~g22665));
assign g27114 = ((~II35297));
assign g11801 = ((~g10988));
assign g5713 = ((~II14163));
assign g22612 = ((~II29194));
assign g30028 = ((~g29567)&(~g29961));
assign g4292 = ((~g2107));
assign g3928 = ((~g157));
assign g28737 = ((~g28428)&(~g27914));
assign g17621 = ((~II23709));
assign g21202 = ((~g19118));
assign II31102 = ((~g22177));
assign g27830 = ((~II36290))|((~II36291));
assign g18217 = ((~g14214));
assign g10627 = (g3678&g5257);
assign II25521 = (g17093)|(g17064)|(g17046);
assign g22570 = ((~II29132));
assign g18508 = ((~g14471));
assign g12453 = ((~II19631));
assign II24595 = ((~g6438))|((~II24594));
assign II34041 = ((~g25566));
assign g11789 = ((~g9480)&(~g9604)&(~g9722));
assign II23518 = ((~g15856));
assign g16411 = (g2593&g12067);
assign g17413 = ((~II23501));
assign g29633 = ((~II39017));
assign g15921 = ((~g12657))|((~g6783));
assign g11926 = (g8169&g8696);
assign g5309 = ((~g2524));
assign g20742 = ((~g20228))|((~g3566));
assign g25037 = ((~g23984))|((~g7195));
assign g12702 = ((~II19794));
assign g19807 = (g1346&g18896);
assign g28696 = ((~II37635));
assign g20434 = ((~g17698));
assign II30029 = ((~g22642));
assign g14040 = (g7691&g12932);
assign g19229 = ((~II25474));
assign g28297 = ((~II37140));
assign g23594 = ((~II30686));
assign II31634 = ((~g23690));
assign II36864 = ((~g27384));
assign g14768 = ((~g12352));
assign g20334 = ((~g17363));
assign g29294 = (g29053&g28900);
assign g30518 = ((~II40134));
assign g20587 = ((~II27086));
assign II23179 = ((~g9488))|((~g13942));
assign g15724 = ((~g12409));
assign g15325 = (g4610&g13197);
assign g13796 = (g7477&g12559);
assign g18853 = ((~g15326));
assign g8899 = (g6945&g1180);
assign II28043 = ((~g19987));
assign g4340 = ((~g343));
assign g25399 = ((~g24787));
assign g10193 = (g3306&g4465);
assign g13936 = ((~g12797));
assign g28258 = ((~II37023));
assign II38142 = ((~g29073));
assign gbuf172 = (g2258);
assign g28810 = ((~II37771));
assign g24886 = ((~II32604));
assign g24246 = (g21982&g11291);
assign g12490 = ((~g8587));
assign g21008 = ((~g19836)&(~g17877));
assign g21480 = (g9795&g20444);
assign II19958 = ((~g8574));
assign g7138 = ((~g2360));
assign g17083 = ((~II23075))|((~II23076));
assign g20997 = ((~g19811)&(~g15487));
assign g23164 = ((~II29945));
assign g21209 = (g20273&g12412);
assign II30607 = ((~g22029));
assign g10361 = (g6448&g4740);
assign g15340 = ((~II21609));
assign g25964 = ((~g22882))|((~g24543));
assign II40721 = ((~g30655));
assign g21987 = ((~g21260)&(~g19541)&(~g19544));
assign II17228 = ((~g7303));
assign g29279 = ((~II38408));
assign g19896 = ((~g16625))|((~g9782));
assign g10829 = ((~g5749));
assign gbuf73 = (g868);
assign g23110 = ((~g17090)&(~g21174));
assign II40766 = ((~g30737));
assign II31478 = ((~g23549));
assign g13515 = (g6044&g12294);
assign g11661 = ((~g9534))|((~g3366));
assign g23710 = ((~II30869))|((~II30870));
assign g10122 = (g3462&g4376);
assign g28880 = (g13946&g28639);
assign II24180 = ((~g9161))|((~II24178));
assign g10189 = ((~II17159));
assign g26121 = ((~II34017));
assign g29613 = ((~g13941)&(~g29257));
assign II25712 = ((~g18048))|((~II25710));
assign g21806 = (g20116)|(g20093)|(g18547)|(g19097);
assign g4329 = ((~g129));
assign II37140 = ((~g28070));
assign g17213 = ((~g4326)&(~g14442));
assign g28075 = ((~II36667))|((~II36668));
assign II36733 = ((~g15055))|((~II36731));
assign g18725 = ((~g13865));
assign g7897 = ((~g3047));
assign g20415 = ((~g17624));
assign g30932 = ((~g30754)&(~g30757));
assign II33608 = ((~g24464));
assign g5327 = ((~g739));
assign II25081 = ((~g14507));
assign g18244 = (g5280&g15741);
assign g28663 = (g27906&g11997);
assign g29885 = ((~g29683));
assign II24586 = ((~g14596))|((~g9488));
assign g13153 = ((~g9199));
assign II30536 = ((~g23081));
assign II24668 = ((~g14559))|((~II24667));
assign II21775 = ((~g13121));
assign g4832 = ((~g1967));
assign II15329 = ((~g3117));
assign II35515 = ((~g26850));
assign II20810 = ((~g13164));
assign g25134 = ((~II32880));
assign g16152 = (g517&g11829);
assign II27128 = ((~g19725));
assign g21716 = ((~g19894));
assign II39407 = ((~g29660));
assign g16312 = (g5870&g11950);
assign g13039 = ((~g9676))|((~g6980));
assign g21674 = ((~g16611)&(~g20025));
assign g24578 = (g1453&g23464);
assign II23807 = ((~g14062))|((~II23806));
assign g8874 = ((~II16138));
assign II38499 = ((~g28772));
assign g12900 = ((~g8941));
assign g26461 = ((~II34421));
assign g13850 = ((~g13386));
assign II33013 = ((~g25119));
assign g30359 = ((~II39892));
assign II35937 = ((~g26822));
assign g26996 = (g23360&g26564);
assign g26495 = ((~II34461));
assign g26775 = (g26099&g22318);
assign g24262 = ((~II31460));
assign g9400 = (g6574&g8076);
assign g15846 = ((~g12611))|((~g6369));
assign g12147 = ((~g8330));
assign g11982 = ((~g11281));
assign g27517 = ((~II35883));
assign g13433 = ((~II20598));
assign g21847 = ((~g13642)&(~g19166));
assign g26119 = ((~g8278))|((~g14657))|((~g25422))|((~g25379));
assign g25549 = ((~II33377));
assign g17855 = (g4839&g15502);
assign II14948 = ((~g2619));
assign g18845 = ((~g15287));
assign II24409 = ((~g14119))|((~II24407));
assign II37854 = ((~g28529));
assign II14808 = ((~g623));
assign g24832 = ((~II32431))|((~II32432));
assign II39071 = ((~g29517));
assign II31751 = ((~g23670));
assign g28949 = (g28630&g9419);
assign g16527 = (g14811&g14849&g16201&g16302);
assign g12466 = ((~g8614));
assign II38101 = ((~g28366));
assign g13999 = ((~g11889));
assign g4380 = ((~g1387));
assign II41123 = ((~g30979));
assign II37044 = ((~g28039));
assign g13117 = ((~g9134));
assign g9955 = (g3722&g4191);
assign g26682 = ((~II34653));
assign g5649 = (g331&g351);
assign g29262 = (g28863&g8965);
assign g24568 = ((~II32112));
assign g9113 = (g3618&g7736);
assign II27314 = ((~g19401));
assign g18999 = ((~II25081));
assign g4220 = ((~g423));
assign g22340 = (g88&g21184);
assign g22684 = ((~II29336));
assign II23153 = ((~g9427))|((~II23152));
assign g8802 = ((~II16006));
assign g8523 = (g6574&g1567);
assign g28459 = (g18074&g27939);
assign g22100 = ((~g21360)&(~g19653));
assign g28053 = ((~II36612));
assign g21522 = (g9857&g20464);
assign g13879 = ((~g11784));
assign g19471 = ((~g18102));
assign g22642 = ((~II29252));
assign g26326 = (g4749&g25585);
assign g22383 = (g1462&g21214);
assign g4951 = ((~g1779));
assign g8503 = (g6314&g270);
assign g4456 = ((~g309));
assign g25986 = ((~II33810));
assign II20431 = ((~g11188))|((~II20429));
assign g11784 = ((~g9463)&(~g9581)&(~g9660));
assign II20688 = ((~g11682));
assign g16880 = ((~g15852)&(~g13056));
assign g25930 = ((~g24978))|((~g5473));
assign g16422 = (g983&g12088);
assign g23244 = ((~II30185));
assign g23844 = ((~II31082));
assign g28287 = ((~II37110));
assign g10631 = ((~g8088));
assign g10182 = (g7488&g4441);
assign g29182 = ((~g28851)&(~g28408));
assign II31586 = ((~g23827));
assign g10437 = (g6678&g4905);
assign g30440 = (g30143&g11095);
assign gbuf125 = (g1786);
assign g24421 = ((~II31937));
assign g30175 = ((~g30020));
assign II24036 = ((~g14016))|((~g9374));
assign g4257 = ((~g1389));
assign II27755 = (g19296&g19478&g19453);
assign g16159 = (g5719&g11835);
assign g10724 = (g3522&g5369);
assign II36120 = ((~g27523));
assign g28373 = (g56&g27969);
assign g15332 = ((~II21601));
assign g30975 = ((~II41099));
assign II24110 = ((~g13963))|((~g9569));
assign g18886 = ((~II24913));
assign g13369 = ((~II20462));
assign g23081 = ((~g17045)&(~g21141));
assign gbuf165 = (g1938);
assign g15245 = (g4474&g13185);
assign II17051 = ((~g3806));
assign II34707 = ((~g26194));
assign g29389 = ((~g29027));
assign II34764 = ((~g26222));
assign g9906 = (g6519&g4130);
assign II38644 = ((~g29299));
assign II21037 = ((~g12486));
assign g10010 = (g6314&g4214);
assign g18341 = ((~g14342));
assign g25445 = ((~g24993));
assign g17091 = (g8004&g15603);
assign g5391 = ((~g2811));
assign g24426 = ((~g23386)&(~g10024));
assign II31814 = ((~g24066));
assign g13702 = (g7802&g12537);
assign g13915 = ((~g8822))|((~g12473))|((~g12463));
assign g4749 = ((~g582));
assign g13320 = (g5685&g11225);
assign g28264 = ((~II37041));
assign II21638 = ((~g11694));
assign g12039 = ((~g11364));
assign g19124 = (g14725&g16656);
assign g29629 = ((~II39005));
assign g18432 = ((~II24459));
assign II30563 = ((~g23111));
assign g16651 = ((~II22694));
assign II36162 = ((~g27385));
assign g8945 = ((~II16247));
assign II30128 = ((~g22828));
assign II38831 = ((~g29324))|((~g15962));
assign II14338 = ((~g2185));
assign II30092 = ((~g22710));
assign g30216 = (g30036&g8921);
assign g21420 = (g9216&g20410);
assign g12079 = ((~g10281)&(~g10361)&(~g10422));
assign g22757 = ((~II29493));
assign II21149 = ((~g13156));
assign g21425 = (g15366&g20416);
assign g26749 = ((~II34854));
assign II29040 = ((~g20693));
assign g30758 = (g30613&g20783);
assign g23642 = ((~II30782));
assign g9441 = (g6314&g8132);
assign g7354 = ((~g1865));
assign g5910 = (g1718&g1705);
assign g15259 = (g4516&g13189);
assign g9422 = ((~II16611));
assign II35539 = ((~g26852));
assign g5786 = (g1718&g1734);
assign g18692 = ((~g14837));
assign g5807 = (g337&g324);
assign g18899 = ((~g15488));
assign g24664 = (g17208&g24134);
assign II32067 = ((~g24174));
assign g29407 = ((~II38606));
assign g13558 = ((~g12657))|((~g3566));
assign g13601 = ((~II20823));
assign g5233 = ((~g620));
assign g26258 = (g4468&g25496);
assign g23229 = ((~II30140));
assign g10059 = (g3566&g4266);
assign g28074 = ((~II36663));
assign g28462 = (g18110&g27946);
assign g26960 = ((~g26597));
assign g30766 = (g30617&g19457&g19431);
assign g24240 = ((~II31426));
assign g28365 = ((~II37260));
assign g26257 = (g4465&g25493);
assign g17548 = ((~II23636));
assign II15986 = ((~g3878));
assign g25802 = ((~II33640));
assign g27522 = ((~II35890));
assign II24054 = ((~g6777))|((~II24053));
assign g30723 = ((~II40459));
assign g11911 = ((~g11170));
assign g16182 = (g7149&g11852);
assign g13401 = ((~g11481)&(~g11332)&(~g7928)&(~g11069));
assign g18503 = ((~g16036)&(~g14464));
assign II36052 = ((~g26954));
assign g3522 = ((~II13194));
assign II24495 = ((~g14048))|((~II24493));
assign II18298 = ((~g6232));
assign II34296 = ((~g25189));
assign g11701 = ((~g9534))|((~g3366));
assign g28282 = ((~II37095));
assign g16938 = (g7858&g15128);
assign g30846 = ((~II40790));
assign g27976 = ((~II36447));
assign g26061 = (g1444&g25315);
assign II21096 = ((~g11749));
assign g23222 = ((~II30119));
assign g26307 = (g4652&g25549);
assign g26762 = ((~II34879));
assign II24679 = ((~g14637))|((~II24677));
assign g21696 = ((~g20487)&(~g7079));
assign g13062 = ((~g9676))|((~g7162));
assign g27140 = ((~g26136));
assign g28310 = ((~II37179));
assign g9108 = (g7015&g7721);
assign g19711 = (g4266&g17531);
assign II35125 = ((~g26096))|((~II35123));
assign g3710 = ((~II13218));
assign g27955 = ((~II36420));
assign II13804 = ((~g2200));
assign g21176 = (g19308&g19295&II27739);
assign g25163 = ((~II32967));
assign g24573 = (g18639&g23129&g23424);
assign II30221 = ((~g22767));
assign g8797 = (g7053&g8009);
assign g23224 = ((~II30125));
assign g27354 = ((~g27112)&(~g26504));
assign g14936 = ((~g12231));
assign g20086 = (g18337&g3170);
assign II24639 = ((~g14390))|((~g15210));
assign g18170 = ((~g15877));
assign II27338 = ((~g19401));
assign g16831 = ((~II22800));
assign g26660 = ((~g25208)&(~g10024));
assign II34449 = ((~g25205));
assign g20346 = ((~g17390));
assign g24488 = ((~g23667)&(~g19740));
assign g17925 = (g4933&g15550);
assign g8576 = (g3722&g2285);
assign II18734 = ((~g9003));
assign g5848 = ((~g2580));
assign II20398 = ((~g10858));
assign g13741 = ((~II20909));
assign g22164 = ((~g21440)&(~g19772));
assign g26986 = (g6438&g26254);
assign g7815 = ((~g2733));
assign g4017 = ((~g427));
assign II17009 = ((~g6945));
assign g28120 = ((~II36789));
assign g19649 = (g4073&g17419);
assign g12291 = ((~g10582)&(~g10624)&(~g10659));
assign g25208 = ((~g24748)&(~g23552));
assign g10281 = (g5438&g4598);
assign g27268 = ((~g26996)&(~g26292));
assign g8539 = (g6574&g1576);
assign g29437 = ((~II38692));
assign g11872 = ((~g9793)&(~g9919)&(~g10055));
assign g10714 = ((~g4495));
assign II34695 = ((~g26167));
assign g12895 = ((~II19952));
assign g8984 = ((~II16300));
assign g11656 = ((~II18842));
assign g22899 = ((~II29690));
assign g16673 = ((~II22715));
assign g12224 = ((~g10469)&(~g10528)&(~g10589));
assign g26082 = (g762&g25771);
assign g28272 = ((~II37065));
assign g5836 = ((~g2297));
assign g23690 = ((~II30854));
assign g13174 = ((~g9351));
assign g20796 = ((~II27385));
assign g19261 = ((~II25533))|((~II25534));
assign g4763 = ((~g731));
assign II23943 = ((~g9293))|((~II23941));
assign g19512 = ((~g17221));
assign gbuf49 = (g325);
assign g24322 = ((~II31640));
assign g14685 = ((~g12245));
assign II18530 = ((~g10888));
assign g24314 = ((~II31616));
assign g10203 = (g6678&g4486);
assign II17681 = ((~g6572));
assign g17019 = ((~II22982))|((~II22983));
assign g12352 = ((~g10673)&(~g10691)&(~g10710));
assign g27626 = ((~g26989))|((~g3306));
assign g21163 = (g19515&g18237&g14431);
assign g15443 = ((~II21705));
assign g13343 = (g5737&g11309);
assign II31847 = ((~g23608));
assign g27324 = ((~g27072)&(~g26424));
assign g19160 = ((~g17446)&(~g15178));
assign g6751 = ((~II14825));
assign II19756 = ((~g10424));
assign g22384 = ((~g21204));
assign II39951 = ((~g30304));
assign g8918 = ((~II16206));
assign II34358 = ((~g25262));
assign II30673 = ((~g22047));
assign II36465 = ((~g27260));
assign g8396 = (g6369&g918);
assign g25152 = ((~II32934));
assign g30749 = ((~II40527));
assign II34713 = ((~g26195));
assign g8031 = ((~II15329));
assign II19560 = ((~g10631));
assign g10430 = (g3338&g4888);
assign II31910 = ((~g23542));
assign g26429 = ((~II34388));
assign II35404 = ((~g26864));
assign II38049 = ((~g28349));
assign II32670 = ((~g23999))|((~II32668));
assign II14925 = ((~g1931));
assign II30735 = ((~g22066));
assign g19299 = ((~g16616));
assign g18756 = ((~g14960));
assign gbuf192 = (g2457);
assign II36609 = ((~g27297));
assign g4561 = ((~g2232));
assign g20108 = (g18543&g3179);
assign II28524 = ((~g21359));
assign g21776 = ((~g20228))|((~g6574));
assign g10011 = (g5438&g4217);
assign g15665 = ((~g12379));
assign g16906 = ((~II22869));
assign II26816 = ((~g17225));
assign g27746 = ((~g27425)&(~g26972));
assign g12021 = ((~g11344));
assign II16700 = ((~g6064));
assign g12246 = ((~g8434));
assign g14885 = ((~g11860));
assign g28898 = (g28619&g9260);
assign g29794 = ((~II39234));
assign g27361 = ((~II35681));
assign g28420 = ((~g16031)&(~g28171));
assign g17526 = (g6421&g16025);
assign g28452 = (g26114&g28166);
assign g29221 = ((~g15305)&(~g28971));
assign g28335 = (g27814&g22343);
assign g16450 = (g5986&g12150);
assign g10393 = (g7195&g1951);
assign g21315 = (g9161&g20313);
assign g12100 = ((~g10307)&(~g10385)&(~g10449));
assign g20021 = (g5369&g18505);
assign gbuf66 = (g549);
assign II19472 = ((~g10683));
assign g29320 = (g29088&g28972);
assign g26245 = ((~II34189));
assign g15604 = (g5162&g13255);
assign g20525 = (g17394&g13849);
assign g9775 = (g6912&g4026);
assign g22958 = ((~g21694));
assign g20365 = ((~g17442));
assign g26675 = ((~g25375)&(~g17176));
assign g21243 = (g19641&g14922&g16712);
assign g17835 = (g4788&g15477);
assign g16575 = ((~g14459));
assign g5193 = ((~g2103));
assign g26186 = (g1372&g25458);
assign II37978 = ((~g28584));
assign g11691 = ((~g9534))|((~g3366));
assign g27016 = (g21983&g26584);
assign g24128 = ((~g22473));
assign g20092 = (g16749&g7603);
assign g21086 = (g20193&g12142);
assign II20577 = ((~g13342));
assign g26581 = ((~g25582));
assign g18223 = (g5260&g15734);
assign g29259 = (g28859&g8925);
assign g10521 = (g7195&g1979);
assign g15808 = ((~g12611))|((~g6519));
assign g4492 = ((~g732));
assign II15922 = ((~g5654));
assign g21140 = (g20095&g14366);
assign g21730 = ((~g20545)&(~g18520));
assign II24206 = ((~g6568))|((~II24205));
assign g6014 = ((~II14475));
assign g19732 = (g660&g18854);
assign II22752 = ((~g14657));
assign g27183 = ((~II35394));
assign II18674 = ((~g9487));
assign II36341 = ((~g27431));
assign II17854 = ((~g6232));
assign II37891 = ((~g28325));
assign g24589 = ((~II32159));
assign g13444 = ((~II20631));
assign II38139 = ((~g29061));
assign g29470 = (g29347&g19530);
assign II35106 = ((~g26675));
assign g23171 = ((~II29966));
assign g22988 = ((~g21404));
assign II30230 = ((~g22796));
assign g29019 = ((~II37978));
assign II35701 = ((~g26867))|((~g26874));
assign II18578 = ((~g8898));
assign g19415 = ((~g16676));
assign g5129 = ((~g2791));
assign II19961 = ((~g10747));
assign g30943 = ((~II41053));
assign II25541 = ((~g18174))|((~II25539));
assign g25996 = ((~II33840));
assign g22589 = ((~II29159));
assign g20752 = ((~g19171)&(~g10238));
assign g29937 = ((~II39411));
assign g20816 = ((~II27405));
assign g15634 = (g5098&g12895);
assign II37047 = ((~g28061));
assign g21065 = ((~g19914)&(~g18169));
assign g10250 = (g7358&g4552);
assign II22842 = ((~g13580));
assign II16811 = ((~g3338));
assign g18992 = ((~II25064));
assign g5148 = ((~g611));
assign g7587 = ((~g2903));
assign g19315 = (g18231)|(g18319);
assign g9585 = ((~II16694));
assign II39902 = ((~g30289));
assign g26809 = ((~g15258)&(~g26270));
assign g5280 = ((~g2790));
assign g27730 = (g27454&g19349);
assign g7855 = ((~II15168))|((~II15169));
assign g17770 = ((~II23845));
assign g26300 = (g4647&g25546);
assign g5179 = ((~g1963));
assign II32444 = ((~g18014))|((~II32443));
assign g30327 = (g30187&g8321);
assign g10408 = (g7303&g2643);
assign II14104 = ((~g331));
assign g24224 = (g22219&g11045);
assign g8677 = ((~II15873));
assign II39369 = ((~g15913))|((~II39367));
assign II20421 = ((~g10808));
assign g26608 = ((~g25669));
assign g24287 = ((~II31535));
assign g25146 = ((~II32916));
assign II13934 = ((~g1060));
assign g27905 = ((~II36358));
assign g13329 = ((~g10337));
assign g13399 = ((~II20505))|((~II20506));
assign g8427 = ((~II15629));
assign g27294 = ((~g27028)&(~g26361));
assign g25387 = ((~g24839));
assign II23584 = ((~g15845));
assign g12690 = ((~g8802));
assign g28677 = ((~II37578));
assign g17031 = (g3410&g10714&g14259);
assign g12121 = ((~g10330)&(~g10406)&(~g10470));
assign g5737 = ((~g1682));
assign g20473 = ((~g18085))|((~g646));
assign g30099 = (g29861&g11287);
assign II40203 = ((~g30380));
assign g5812 = ((~g915));
assign g29243 = (g9857&g28829);
assign g14286 = ((~g12048));
assign g23778 = (g22954&g9531);
assign g24146 = ((~g22509));
assign g13867 = ((~g11773));
assign g6231 = ((~II14712));
assign g19105 = ((~II25294));
assign g10494 = (g6643&g608);
assign g26959 = ((~II35146));
assign II40898 = ((~g30832));
assign g25226 = ((~g24774)&(~g23584));
assign g7534 = ((~g1832));
assign g7529 = ((~g465));
assign g28400 = ((~g27886)&(~g22344));
assign g3678 = ((~II13215));
assign g22191 = ((~g21517)&(~g19850));
assign g11981 = ((~g10117)&(~g10207)&(~g10294));
assign g12125 = ((~II19307));
assign g22775 = ((~II29539));
assign g24068 = ((~II31290));
assign II36258 = ((~g15859))|((~II36256));
assign g29346 = (g29087&g29077);
assign g20711 = ((~II27300));
assign g26571 = ((~g25554));
assign g17024 = ((~II22999))|((~II23000));
assign g5207 = ((~g2649));
assign g28187 = ((~g27543));
assign II28994 = ((~g21715));
assign II26538 = (g18319)|(g18231)|(g18147);
assign g16803 = ((~g15593)&(~g12908));
assign II17969 = ((~g5880));
assign g9367 = (g6232&g8062);
assign g13360 = (g5766&g11373);
assign g26283 = ((~g25954)&(~g24486));
assign g24770 = ((~g16119)&(~g24217));
assign g12801 = ((~II19862));
assign II13655 = ((~g2175));
assign g19869 = (g679&g18926);
assign II23475 = ((~g15821));
assign g5164 = ((~g1405));
assign g17149 = (g7694&g14115);
assign II33188 = ((~g24814));
assign g25125 = ((~g23510)&(~g22340));
assign g18650 = (g14976&g16201&g16302);
assign g29501 = ((~II38827));
assign g30284 = ((~g16444)&(~g29980));
assign II40781 = ((~g30808));
assign g10377 = (g6945&g4780);
assign g5050 = ((~g1269));
assign g16082 = ((~g10952)&(~g6140)&(~g12487));
assign g22907 = ((~g21711));
assign g22876 = ((~g21238))|((~g83));
assign g26816 = ((~g15351)&(~g26312));
assign II37358 = ((~g27811))|((~II37356));
assign II39050 = ((~g29515));
assign g11538 = ((~II18590));
assign g11509 = ((~II18503));
assign g27783 = (g5819&g27373);
assign g17738 = ((~II23817));
assign g5304 = ((~g1991));
assign g30367 = (g30207&g8460);
assign g10214 = ((~II17184));
assign II34797 = ((~g26208));
assign g26618 = ((~II34579));
assign II32286 = ((~g23953))|((~II32284));
assign g8381 = ((~g8182))|((~g8120))|((~g8044))|((~g7989));
assign II18214 = ((~g3254));
assign g14280 = ((~g12044));
assign g16611 = ((~g15962)&(~g15942)&(~g15923));
assign g30477 = (g30183&g11321);
assign g28919 = (g14107&g28644);
assign g12931 = ((~g8965));
assign II32567 = ((~g18131))|((~g24082));
assign II34077 = ((~g25954));
assign g17226 = ((~g16010)&(~g16017));
assign g19054 = ((~II25225));
assign g24331 = ((~II31667));
assign g28362 = ((~g15730)&(~g28105));
assign g18371 = ((~II24394));
assign II37822 = ((~g28384))|((~g28386));
assign II26708 = (g18699&g18728&g16201);
assign g11160 = ((~II18076));
assign g9737 = ((~g5834));
assign II34080 = ((~g25539));
assign g20248 = (g18656&g14837&g16293);
assign g11994 = ((~g11300));
assign g4848 = ((~g2257));
assign g23782 = ((~II30988));
assign g12836 = ((~g8417)&(~g8458)&(~g8481));
assign g24207 = ((~g16967)&(~g22229));
assign g29480 = (g21461&g29282);
assign g6974 = ((~g1151));
assign II25923 = ((~g18526))|((~II25921));
assign g7664 = ((~g2387));
assign g28111 = (g27617&g10263);
assign g27482 = ((~g26906)&(~g24637));
assign g28580 = ((~II37497));
assign g25752 = ((~II33583));
assign g26012 = ((~II33888));
assign g28309 = ((~II37176));
assign II39068 = ((~g29516));
assign II15532 = ((~g3410));
assign g21586 = ((~II28115));
assign II35049 = ((~g26530));
assign g24372 = ((~II31790));
assign g11330 = ((~II18281))|((~II18282));
assign g25096 = ((~g23979))|((~g1365));
assign g23550 = (g8132&g22409);
assign II18512 = ((~g9309));
assign g10238 = (g3710&g7358);
assign g20921 = ((~g19697)&(~g17576));
assign II30928 = ((~g22128));
assign g25288 = ((~g24938)&(~g18256));
assign g16985 = ((~II22918))|((~II22919));
assign g14148 = ((~g12912));
assign g26742 = ((~II34833));
assign II33580 = ((~g25051));
assign g8937 = ((~II16231));
assign g11908 = ((~g11160));
assign g10295 = (g3462&g4641);
assign g4548 = ((~g1810));
assign II23083 = ((~g9310))|((~II23082));
assign g8012 = ((~II15304));
assign II37107 = ((~g28043));
assign g27386 = ((~g27143));
assign g27566 = ((~II35975))|((~II35976));
assign g8756 = ((~II15946));
assign g13025 = ((~g10810));
assign g23857 = (g14263&g23056);
assign g30715 = ((~II40435));
assign g15385 = ((~II21647));
assign g21067 = (g20193&g12030);
assign g21723 = (g3554&g20534);
assign g22283 = ((~g20729));
assign g22461 = ((~II29007));
assign g10708 = ((~g3710))|((~g7358));
assign g5656 = ((~g987));
assign g24052 = ((~g22812))|((~g14171));
assign g29574 = ((~g28712)&(~g29180));
assign II38872 = ((~g29182));
assign g22319 = ((~g21228));
assign g13195 = ((~g9524));
assign II15806 = ((~g5550));
assign g8000 = ((~g853));
assign g27997 = ((~g16456)&(~g27242));
assign II15850 = ((~g5627));
assign g21558 = ((~II28090));
assign g30104 = (g29853&g11361);
assign g24582 = ((~II32140));
assign g21822 = (g16778&g19681&g14936);
assign g28704 = ((~II37659));
assign g3806 = ((~II13232));
assign II23143 = ((~g9407))|((~II23142));
assign g11795 = ((~g10977));
assign g21467 = ((~g20506)&(~g13355));
assign g28044 = ((~II36585));
assign II38250 = ((~g28941));
assign g7338 = ((~g3002));
assign g15553 = ((~II21809));
assign g23551 = (g8135&g22412);
assign g26737 = ((~II34818));
assign g20928 = ((~g19921));
assign II25856 = ((~g1453))|((~II25855));
assign g21107 = (g19444&g17893&g14079);
assign II34946 = ((~g26534));
assign g16016 = (g5601&g11740);
assign II14763 = ((~g405));
assign g7229 = ((~II14934));
assign II39631 = ((~g30084));
assign g5551 = ((~g514));
assign g22694 = ((~II29354));
assign g27297 = ((~g27031)&(~g26365));
assign g15262 = ((~g12204));
assign g23277 = ((~II30284));
assign g19209 = (g18079)|(g18346);
assign g12430 = ((~g10905));
assign g24523 = ((~g23842)&(~g22714));
assign g21871 = ((~g18458))|((~g19225))|((~g19232));
assign g17718 = (g4451&g16064);
assign g14183 = ((~II21108));
assign g25412 = ((~g24791));
assign g29112 = ((~g28661)&(~g17100));
assign g14795 = ((~II21318));
assign g5939 = ((~g1627));
assign II13896 = ((~g343));
assign g4552 = ((~g2086));
assign g26157 = (g21825&g25630);
assign gbuf187 = (g2432);
assign g23872 = ((~II31130));
assign g29300 = (g29072&g28925);
assign g24341 = ((~II31697));
assign II36960 = ((~g28011));
assign g25588 = ((~II33411));
assign g26645 = ((~g25808));
assign g26508 = ((~g25312));
assign II22524 = ((~g13673));
assign g24754 = (g15540&g24107);
assign II32547 = ((~g17903))|((~II32546));
assign g5057 = ((~g1291));
assign g7879 = ((~g3065));
assign g8517 = (g6232&g204);
assign g26719 = ((~II34764));
assign g30308 = ((~II39767));
assign g29686 = ((~g29566)&(~g29342));
assign g29097 = ((~g28335)&(~g28336));
assign g22887 = ((~II29687));
assign g26498 = ((~g25372))|((~g1439));
assign g24880 = ((~II32587))|((~II32588));
assign II29351 = ((~g20963));
assign g20447 = ((~g17764));
assign g23359 = ((~g22216)&(~g22907));
assign II26667 = (g14922&g18765&g13724);
assign g20971 = ((~II27516));
assign g23557 = ((~II30617));
assign II32871 = ((~g24518));
assign g20570 = ((~II27035));
assign II39638 = ((~g30056));
assign g20241 = (g13764&g13819&II26667);
assign II30284 = ((~g22662));
assign g14431 = ((~g12121));
assign g30504 = (g30183&g11462);
assign II37804 = ((~g28636));
assign g30072 = ((~g29910)&(~g8947));
assign g19902 = (g14201&g18368&II26348);
assign g6519 = ((~II14778));
assign II21364 = ((~g13028));
assign g6100 = ((~II14615));
assign g23588 = ((~II30676));
assign II28155 = (g14033&g14472&g14107);
assign II27391 = ((~g19420));
assign g25378 = ((~g24877));
assign g10329 = (g3774&g4721);
assign g21118 = ((~g20091)&(~g20113)&(~g20136));
assign g24432 = (g14642&g15904&g24115);
assign g21123 = (g19970&g19982);
assign II34505 = ((~g25450));
assign g11865 = ((~g9781)&(~g9909)&(~g10045));
assign g19941 = (g2760&g18974);
assign g26657 = ((~g25862));
assign g5622 = ((~g3176));
assign g17051 = ((~g14657)&(~g15880)&(~g14630));
assign g19796 = (g2727&g18881);
assign II15651 = ((~g3722));
assign g18369 = ((~II24381))|((~II24382));
assign II28162 = (g18142&g18526&g18226);
assign g21878 = ((~g16964)&(~g19228));
assign g22247 = ((~g21695)&(~g20001));
assign II28174 = ((~g20025));
assign II26396 = (g18585&g14234&g14332);
assign II23712 = ((~g15872));
assign g5775 = ((~g1481));
assign g24405 = ((~II31889));
assign g24656 = ((~g23715)&(~g22624));
assign g16507 = ((~g14186));
assign g14641 = ((~g11823));
assign g11271 = ((~II18217));
assign II14618 = ((~g2459));
assign II34124 = ((~g25225));
assign II36426 = ((~g27584));
assign g28863 = ((~g28417));
assign II14605 = ((~g468));
assign II17774 = ((~g8107));
assign g24904 = ((~II32646))|((~II32647));
assign g27548 = ((~II35940));
assign g29395 = ((~g29054));
assign II39800 = ((~g30309));
assign II40128 = ((~g30479));
assign g23953 = ((~g22812))|((~g14525));
assign g13166 = ((~g9290));
assign g21455 = (g15366&g20436);
assign g11410 = ((~II18369))|((~II18370));
assign g25233 = ((~g24788)&(~g23604));
assign g7712 = ((~g1089));
assign g29142 = ((~II38169));
assign g4211 = ((~g159));
assign g22080 = ((~g21344)&(~g19624));
assign II30725 = ((~g22064));
assign II29375 = ((~g20969));
assign g25013 = ((~g23923))|((~g6643));
assign II18452 = ((~g10930));
assign II37295 = ((~g27827))|((~g27814));
assign g11737 = ((~g10809));
assign g8931 = ((~II16221));
assign g26730 = ((~II34797));
assign g28163 = ((~g27437));
assign II22918 = ((~g15096))|((~II22917));
assign g10678 = (g6912&g5327);
assign g15877 = ((~g13374))|((~g12392));
assign g12370 = ((~II19530));
assign II15543 = ((~g3410));
assign g25859 = ((~II33703));
assign g29361 = ((~g28877));
assign g18796 = ((~g15080));
assign II38474 = ((~g28759));
assign g26635 = ((~g25758));
assign g29755 = ((~g16229)&(~g29610));
assign II14577 = ((~g1836));
assign g29609 = ((~g13900)&(~g29252));
assign II38496 = ((~g28771));
assign g28174 = ((~g27489));
assign g16264 = (g5822&g11909);
assign II27822 = ((~g19865));
assign g25400 = ((~g24712));
assign g29317 = ((~II38480));
assign II16015 = ((~g6056));
assign II32961 = ((~g24851));
assign II31499 = ((~g23588));
assign II19208 = ((~g10424));
assign g26613 = ((~g25685));
assign II26357 = (g18469&g18573&g18314);
assign g30285 = ((~g16447)&(~g29981));
assign g5953 = ((~g97));
assign II34983 = ((~g26569));
assign g27033 = (g23364&g26604);
assign g27023 = (g23349&g26591);
assign II29310 = ((~g20947));
assign II40618 = ((~g30566));
assign g13184 = ((~g9419));
assign g27707 = ((~II36132));
assign II25809 = ((~g767))|((~g17993));
assign g14028 = ((~g11905));
assign g28223 = ((~II36918));
assign g10510 = (g6751&g1291);
assign g24443 = ((~g23644))|((~g3306));
assign II18277 = ((~g7391));
assign g21932 = ((~II28447));
assign g24412 = ((~II31910));
assign g17255 = ((~II23341));
assign g5604 = ((~g3167));
assign g27962 = ((~g16394)&(~g27679));
assign g13463 = ((~II20688));
assign g23860 = (g22962&g9790);
assign g23160 = ((~II29933));
assign II26676 = (g18708&g18735&g16266);
assign g20116 = (g16142&g13677&g13706&II26558);
assign II38352 = ((~g29110));
assign g30293 = ((~g13480)&(~g29989));
assign g20085 = (g18170&g3164);
assign g16483 = ((~II22551));
assign g19190 = ((~II25415));
assign II32988 = ((~g24589));
assign g5895 = ((~g255));
assign g25732 = ((~II33561));
assign g25513 = (g24487&g17664);
assign g24472 = ((~g24014))|((~g3806));
assign g15094 = (g7872&g12604);
assign II39089 = ((~g29495));
assign g17151 = ((~g14753)&(~g15971)&(~g14711));
assign g22999 = ((~g21085)&(~g19241));
assign g12504 = ((~g8643));
assign II26500 = (g18465&g18389&g18313);
assign II37912 = ((~g28584));
assign g17882 = ((~g13946));
assign II27203 = ((~g20491));
assign g27814 = ((~g6087)&(~g27632)&(~g25322));
assign g18414 = ((~g15718));
assign g13499 = (g6034&g12252);
assign g28567 = (g26512)|(g27751);
assign g29281 = ((~II38412));
assign g13218 = ((~g9767));
assign g28340 = (g28088&g19519);
assign g23900 = (g22980&g9965);
assign g27759 = ((~g27495)&(~g27052));
assign g25052 = ((~g24014))|((~g7391));
assign g11880 = (g6294&g8678);
assign g5408 = ((~II13940));
assign II38483 = ((~g28990));
assign g11007 = ((~II17916));
assign g8564 = (g3722&g2267);
assign g16107 = (g5666&g11801);
assign II26545 = ((~g16823));
assign g24558 = ((~g23917)&(~g22804));
assign g19787 = (g18038&g16062);
assign g10650 = (g6678&g5293);
assign II22763 = ((~g14753));
assign g22139 = ((~g21397)&(~g19719));
assign g19970 = (g18354&g18276&II26416);
assign II23217 = ((~g9613))|((~g13903));
assign gbuf210 = (g2602);
assign II30829 = ((~g22098));
assign II28485 = ((~g21426));
assign gbuf83 = (g973);
assign II33526 = ((~g24457));
assign g29303 = ((~g28716)&(~g19112));
assign II19557 = ((~g10606));
assign g4427 = ((~g2236));
assign g26396 = (g5027&g25700);
assign g19842 = (g14525&g13922&II26282);
assign g24004 = ((~g4809)&(~g13582)&(~g23042));
assign II36867 = ((~g27786));
assign g30647 = ((~g16251)&(~g30447));
assign g13421 = ((~II20562));
assign II17945 = ((~g5668));
assign g19204 = (g18556)|(g18115);
assign II13913 = ((~g373));
assign II36141 = ((~g27559));
assign g10044 = (g6369&g4243);
assign g5662 = ((~g2589));
assign II35476 = ((~g27163));
assign II35923 = ((~g26820));
assign g5389 = ((~g3040));
assign g12851 = ((~g8888));
assign g24604 = (g1457&g23908);
assign II29408 = ((~g20980));
assign g30131 = (g30059&g20749);
assign g25530 = ((~II33358));
assign g16702 = ((~II22730));
assign g24551 = ((~II32085));
assign g23233 = ((~II30152));
assign II34063 = ((~g25209));
assign II19488 = ((~g10653));
assign g29881 = ((~g29682));
assign g29555 = (g29224&g29387);
assign II23208 = ((~g9595))|((~II23207));
assign g12008 = ((~g10183)&(~g10270)&(~g10351));
assign g30728 = (g30605&g22252);
assign g24280 = ((~II31514));
assign g29398 = ((~g29069));
assign g28416 = (g7823&g27889);
assign g25139 = ((~II32895));
assign II37920 = ((~g28501));
assign g21414 = (g15118&g20406);
assign g16187 = (g5754&g11857);
assign g6212 = ((~g1378));
assign g5951 = ((~II14413));
assign g12142 = ((~II19321));
assign g9112 = (g3462&g7733);
assign g9306 = ((~II16541));
assign g4507 = ((~II13501));
assign II22683 = ((~g14725));
assign II33801 = ((~g25327));
assign g25073 = ((~g24014))|((~g7391));
assign II18108 = ((~g7855))|((~II18106));
assign g21023 = ((~g19855)&(~g15573));
assign g30263 = ((~g16344)&(~g30097));
assign g9419 = ((~II16608));
assign g8654 = (g3806&g7484);
assign g13095 = ((~g10839));
assign g10166 = (g7230&g4415);
assign g5746 = ((~g2375));
assign II23345 = ((~g15723));
assign g23771 = (g22720&g20455);
assign g13427 = ((~II20580));
assign g18720 = ((~g14895));
assign g29974 = ((~II39460));
assign II30185 = ((~g22658));
assign II38999 = ((~g29496));
assign g23910 = (g22971&g10067);
assign g27775 = (g5790&g27506);
assign II38716 = ((~g29230));
assign II21497 = ((~g11674));
assign II20604 = ((~g12440));
assign g28681 = ((~II37590));
assign g27413 = ((~g27038))|((~g7015));
assign g25443 = ((~II33268));
assign g26168 = ((~g25953)&(~g16212));
assign g3237 = ((~II13107));
assign g12429 = (g8101&g9044);
assign g16014 = ((~g12695));
assign g19026 = ((~II25141));
assign g9123 = (g3774&g7766);
assign II29690 = ((~g21080));
assign g19722 = (g2714&g18849);
assign II37330 = ((~g28194));
assign gbuf24 = (g180);
assign g26407 = ((~II34369));
assign g26295 = ((~g25977)&(~g13385));
assign g11382 = ((~II18338));
assign g10617 = ((~g8083));
assign g8665 = ((~II15859));
assign g29663 = ((~g29518)&(~g29284));
assign g10548 = (g3306&g5142);
assign g5504 = ((~g3086));
assign g4725 = ((~g2775));
assign g23726 = (g21825&g22843);
assign g25426 = ((~g24183)&(~g24616));
assign g5627 = ((~g125));
assign g24704 = ((~g23509));
assign g24254 = (g19454)|(g22403);
assign g18655 = (g14936&g15161&g16325&g13840);
assign g25776 = ((~II33611));
assign g20388 = ((~g17523));
assign g26386 = (g4994&g25685);
assign g15127 = (g4250&g13170);
assign II16544 = ((~g6054));
assign g23432 = (g21631&g22476);
assign g7766 = ((~g2477));
assign g15353 = ((~g12256));
assign II13152 = ((~g48));
assign g10107 = (g5438&g438);
assign II27491 = ((~g20314));
assign g26144 = ((~g23803))|((~g25402));
assign g8502 = (g3254&g264);
assign g12955 = (g9822)|(g3710);
assign g23531 = ((~II30575));
assign g18810 = ((~g15133));
assign II21523 = ((~g13069));
assign g23158 = ((~II29927));
assign II25092 = ((~g14423));
assign g22177 = ((~g21476)&(~g19806));
assign g10331 = ((~g5366));
assign g13418 = ((~II20553));
assign II22702 = ((~g14737));
assign II26320 = (g18374&g18509&g18207);
assign g17433 = ((~II23521));
assign g11763 = ((~g10918));
assign g19227 = (g18478)|(g18531);
assign II19321 = ((~g10549));
assign g10112 = (g3366&g4348);
assign II23863 = ((~g15151));
assign II33374 = ((~g25031));
assign g10866 = ((~g5849));
assign II36936 = ((~g28072));
assign g24530 = ((~g23857)&(~g22732));
assign II36367 = ((~g27678));
assign g4282 = ((~g1798));
assign II21936 = ((~g13128));
assign g30336 = ((~II39843));
assign g19288 = ((~g14685))|((~g8580))|((~g17057));
assign II23588 = ((~g14885));
assign II33825 = ((~g25462));
assign g7956 = ((~II15262));
assign g30773 = ((~II40581));
assign g9807 = (g6783&g4058);
assign g26415 = (g5081&g25738);
assign g19747 = (g4395&g17607);
assign g20341 = ((~g17375));
assign II27426 = ((~g19457));
assign g16324 = (g5879&g11960);
assign g21598 = ((~g19309));
assign g28983 = ((~II37950));
assign II29212 = ((~g20912));
assign II26134 = ((~g18201));
assign g7460 = ((~g1471));
assign II14599 = ((~g2444));
assign g5819 = ((~g1430));
assign g26798 = ((~g26055)&(~g18407));
assign g24512 = ((~g23795)&(~g22679));
assign g29764 = ((~g16462)&(~g29464));
assign g17796 = (g4728&g15446);
assign II24923 = ((~g14849));
assign g9080 = (g5473&g7658);
assign g8059 = ((~g148));
assign II27002 = ((~g19147));
assign II21446 = ((~g13029));
assign g24111 = ((~g22440));
assign II16469 = ((~g7936));
assign II36696 = ((~g27321));
assign g5098 = ((~g2111));
assign II25554 = (g17131)|(g17099)|(g17080);
assign II29566 = ((~g21039));
assign II15481 = ((~g3248));
assign g18539 = ((~II24608));
assign g8255 = ((~g3072));
assign g26221 = ((~II34153));
assign g11947 = ((~g10061)&(~g10152)&(~g10223));
assign g13147 = ((~g8278))|((~g3306));
assign g10968 = ((~II17863));
assign g30011 = ((~g29522)&(~g29944));
assign II38258 = ((~g28963));
assign II23670 = ((~g15912));
assign g19444 = ((~g17985));
assign g23211 = ((~II30086));
assign g27330 = ((~g27082)&(~g26441));
assign II33219 = ((~g24849));
assign g19593 = (g8239&g17336);
assign g26756 = (g26113&g22240);
assign g28292 = ((~II37125));
assign g26690 = ((~II34677));
assign g18894 = ((~g15471));
assign g13492 = (g2371&g12222);
assign g6777 = ((~g1346));
assign g16062 = ((~g12801));
assign II23027 = ((~g15366))|((~g14221));
assign g15700 = (g5279&g13284);
assign II18085 = ((~g5611));
assign g29511 = ((~II38863));
assign g19352 = ((~II25751))|((~II25752));
assign g17182 = (g8084&g15792);
assign g8587 = ((~g6418));
assign g14321 = ((~g12062));
assign g23562 = ((~II30626));
assign g20103 = (g18332&g18257&II26541);
assign II37125 = ((~g28090));
assign g12650 = (g6149&g9290);
assign g13901 = ((~g11810));
assign II25872 = ((~g17183));
assign g25099 = ((~g23440)&(~g22224));
assign g25947 = ((~g24554)&(~g24563));
assign II32295 = ((~g18014))|((~g23968));
assign g18957 = ((~g13884)&(~g12307));
assign g12421 = ((~II19569));
assign g15429 = ((~II21691));
assign g18914 = ((~g15547));
assign g11327 = ((~II18277));
assign g26701 = ((~II34710));
assign g28732 = ((~g14894)&(~g28426));
assign g22699 = (g7338&g21883);
assign II19552 = ((~g8430));
assign g15458 = ((~g12312));
assign g30964 = ((~g30961));
assign g22590 = ((~II29162));
assign g20336 = ((~g17369));
assign g28206 = ((~II36867));
assign II31739 = ((~g23668));
assign g27337 = ((~g27089)&(~g26456));
assign g7475 = ((~g493));
assign g15561 = (g5087&g13239);
assign g15888 = ((~g12611))|((~g6519));
assign g19131 = (g14753&g16673);
assign II32439 = ((~g23392));
assign g28357 = ((~g15681)&(~g28087));
assign g26030 = (g25429&g22304);
assign g28488 = ((~g26755)&(~g27719));
assign g10226 = (g3618&g1804);
assign g18929 = ((~g15609));
assign II27240 = ((~g19335));
assign g28707 = (g12436&g28379);
assign II18166 = ((~g5778));
assign II18157 = ((~g3566));
assign g26935 = ((~g26327));
assign g8273 = ((~II15487));
assign II30991 = ((~g22146));
assign g21521 = (g9941&g20463);
assign g4324 = ((~g2867));
assign g6712 = ((~II14816));
assign g28747 = ((~g28434)&(~g27923));
assign g8912 = ((~II16200));
assign g9056 = (g6945&g1253);
assign g13103 = ((~g9676))|((~g7162));
assign g30314 = ((~II39785));
assign g24466 = ((~g23984))|((~g3650));
assign II39773 = ((~g30064));
assign g29692 = ((~II39130));
assign g23207 = ((~II30074));
assign II27131 = ((~g19798));
assign g10644 = (g7426&g5286);
assign g29416 = ((~II38629));
assign II29001 = ((~g20658));
assign g18634 = ((~g16278));
assign g27743 = ((~g25384))|((~g27436));
assign g23603 = ((~II30707));
assign II17727 = ((~g7013));
assign g12268 = ((~g10529)&(~g10590)&(~g10629));
assign g19533 = ((~g16832));
assign II24437 = ((~g14153))|((~II24436));
assign gbuf96 = (g1082);
assign II38018 = ((~g28342));
assign II38713 = ((~g29410));
assign g22664 = ((~II29294));
assign g21376 = ((~II27917));
assign II39534 = ((~g29917))|((~II39532));
assign g4929 = ((~g1285));
assign g20137 = (g18070&g9226);
assign g19880 = (g2046&g18934);
assign II37161 = ((~g28120));
assign g24303 = ((~II31583));
assign g11935 = ((~g10014)&(~g10106)&(~g10196));
assign g16813 = ((~II22783));
assign g13528 = ((~g12565))|((~g3254));
assign g24461 = ((~g23984))|((~g3650));
assign g22936 = ((~g21255))|((~g1457));
assign g9096 = (g6713&g7685);
assign g16212 = (g5609&g13252);
assign g25160 = ((~II32958));
assign g13072 = ((~g9534))|((~g6912));
assign g7614 = ((~g2543));
assign g16283 = (g5836&g11919);
assign g27122 = ((~g26410))|((~g7015));
assign g26638 = ((~g25776));
assign gbuf12 = (g2836);
assign g13292 = ((~II20351));
assign II14535 = ((~g2546));
assign g22005 = ((~g21540))|((~g21572));
assign g5110 = ((~g2473));
assign II23817 = ((~g13557));
assign II35355 = ((~g26130));
assign g29523 = (g28737&g29364);
assign g15439 = ((~g12299));
assign g24408 = ((~II31898));
assign g9076 = (g5438&g7646);
assign gbuf197 = (g2406);
assign II20523 = ((~g13317));
assign g12059 = ((~II19240));
assign g17117 = (g7906&g15665);
assign II30137 = ((~g22591));
assign g9464 = (g6369&g8147);
assign g23743 = (g6777&g23015);
assign g29411 = (g29090&g21932);
assign II24894 = ((~g14797));
assign g24103 = ((~g22397));
assign g22700 = (g7146&g21558);
assign II14888 = ((~g1925));
assign g10986 = ((~g6014));
assign g25793 = ((~II33630));
assign II18197 = ((~g7896))|((~g7876));
assign g13892 = (g7616&g12815);
assign g19540 = (g16884&g16697&g14797);
assign g9391 = ((~g5867));
assign g5593 = ((~g789));
assign g27761 = ((~g27516)&(~g27079));
assign II19342 = ((~g10574));
assign II23845 = ((~g16174));
assign g26672 = ((~g25365)&(~g17172));
assign II28152 = ((~g20025));
assign g6305 = ((~g2760));
assign g29751 = ((~g6104)&(~g29583)&(~g25352));
assign g26067 = (g25946&g21125);
assign g17436 = ((~II23524));
assign g4104 = ((~g163));
assign g30802 = ((~II40658));
assign g5736 = ((~g1594));
assign g22724 = ((~II29418));
assign g22397 = ((~g14618))|((~g21204))|((~g10754));
assign II16221 = ((~g5412));
assign g23146 = ((~g21825));
assign II30107 = ((~g22735));
assign g30614 = ((~g6119)&(~g30412)&(~g25403));
assign g26586 = ((~g25596));
assign g10351 = (g3834&g4725);
assign g30863 = ((~II40841));
assign II35153 = ((~g26677));
assign g10817 = ((~II17662));
assign g21954 = ((~II28488));
assign g16043 = ((~g12769));
assign g9607 = ((~II16711));
assign g24370 = ((~II31784));
assign g19212 = (g18290)|(g18497);
assign II21580 = ((~g13053));
assign g10076 = (g3722&g4295);
assign g21309 = (g9310&g20304);
assign g19930 = (g2760&g18966);
assign g4683 = ((~II13575));
assign g5341 = ((~g2685));
assign g24591 = (g83&g23853);
assign g16385 = (g5714&g13336);
assign II26476 = ((~g17111));
assign g4147 = ((~g1386));
assign g18865 = ((~g15385));
assign g23765 = ((~II30959));
assign g22608 = ((~g20842))|((~g20885));
assign g8009 = ((~g1869));
assign g23923 = ((~II31195));
assign g7721 = ((~g1785));
assign II18629 = ((~g8811));
assign g22519 = ((~II29067));
assign g15197 = (g4379&g13179);
assign g16442 = ((~g12565))|((~g3254));
assign g27161 = ((~II35360));
assign g28449 = ((~g27727)&(~g26780));
assign g24882 = (g1352&g23832);
assign g19811 = (g18014&g16091);
assign g14613 = ((~g12272));
assign g28157 = ((~g13902)&(~g27370));
assign g30912 = ((~II40988));
assign g21886 = ((~g19915));
assign II36563 = ((~g27286));
assign g5858 = ((~g771));
assign II33361 = ((~g25013));
assign g18036 = (g5092&g15628);
assign g21735 = (g3866&g20536);
assign II25692 = ((~g17741))|((~II25690));
assign g15221 = ((~g12166));
assign g23100 = (g21821)|(g21817)|(g21856);
assign g23591 = (g4012&g22480);
assign g30686 = ((~g16461)&(~g30340));
assign g12907 = ((~g8949));
assign g11490 = ((~g8276));
assign g13348 = ((~II20430))|((~II20431));
assign g11777 = ((~g10946));
assign II36246 = ((~g27674));
assign II16252 = ((~g6134));
assign g10629 = (g3774&g5263);
assign g15115 = ((~II21435));
assign g9857 = ((~g5793));
assign g4994 = ((~g2421));
assign g23308 = ((~II30377));
assign g19418 = ((~g17162));
assign g30979 = ((~II41111));
assign II38154 = ((~g29089));
assign g23891 = (g14385&g23074);
assign II37386 = ((~g28194));
assign g19383 = ((~g16659));
assign II37650 = ((~g28347));
assign g30786 = ((~g30625)&(~g22387));
assign g22647 = ((~II29259));
assign g23730 = ((~II30914));
assign g27166 = ((~II35369));
assign g21041 = ((~g19881)&(~g18037));
assign II25742 = ((~g17842))|((~II25740));
assign g24687 = ((~g23493));
assign II18217 = ((~g6314));
assign g18903 = ((~g15510));
assign II13366 = ((~g2851));
assign g20007 = ((~g18639));
assign g26820 = ((~g15423)&(~g26346));
assign g24675 = ((~g23769)&(~g22660));
assign g1942 = ((~II13095));
assign g27854 = ((~g27632)&(~g1218));
assign II21531 = ((~g11683));
assign II26985 = ((~g16943));
assign g20598 = ((~II27119));
assign g29536 = (g29207&g29375);
assign g30115 = (g29873&g11450);
assign g5762 = ((~g906));
assign g18668 = (g15161&g16325&g16404);
assign II22557 = ((~g14775));
assign g14570 = ((~g12232));
assign II36714 = ((~g27326));
assign II17156 = (g6898&g2998&g6901&g3002);
assign II18560 = ((~g8844));
assign g30373 = ((~II39926));
assign g8808 = ((~II16012));
assign II36653 = ((~g27310));
assign g24211 = (g22014&g10969);
assign g10800 = ((~II17645));
assign g5873 = (g1712&g1777);
assign g10921 = ((~II17804));
assign g21093 = ((~g19075));
assign g24115 = ((~g22381));
assign g25241 = ((~g24799)&(~g23623));
assign g25870 = ((~g4456)&(~g25078)&(~g18429)&(~g16075));
assign II30757 = ((~g22075));
assign g9132 = (g5512&g7792);
assign g8824 = ((~II16044));
assign g25085 = ((~g23432)&(~g22208));
assign II18491 = ((~g8891));
assign g25981 = (g24819&g13858);
assign II18229 = ((~g3410));
assign II28521 = ((~g21824));
assign g4254 = ((~g1384));
assign g11966 = (g8090&g8708);
assign g13787 = (g7967&g11923);
assign II36354 = ((~g27662));
assign g23660 = ((~II30791))|((~II30792));
assign g15922 = ((~g12657))|((~g6574));
assign II21998 = ((~g11729));
assign II27077 = ((~g19259));
assign g20577 = ((~II27056));
assign II17734 = ((~g7138));
assign II25456 = ((~g18883));
assign g28713 = (g28410&g22290);
assign II37514 = ((~g27771));
assign g7718 = ((~g1699));
assign g9965 = ((~II16961));
assign g16996 = ((~II22953))|((~II22954));
assign g20219 = (g16371&g13825&II26654);
assign g10659 = (g3650&g5301);
assign II40119 = ((~g30435));
assign g14959 = ((~g11976));
assign g28006 = ((~II36499));
assign g13646 = (g7772&g12505);
assign g17357 = ((~II23445));
assign II13910 = ((~g361));
assign g9958 = ((~II16954));
assign g18278 = ((~II24285));
assign g29185 = ((~g28853)&(~g28412));
assign II32511 = ((~g24070))|((~II32509));
assign g23720 = ((~II30894));
assign g16010 = (g7639&g11736);
assign g8475 = ((~II15677));
assign g22376 = ((~II28928));
assign g24548 = ((~g15640)&(~g23915));
assign II31031 = ((~g22576));
assign g17627 = ((~II23715));
assign II13901 = ((~g346));
assign g14027 = ((~g10749))|((~g12490));
assign g16251 = (g5812&g11898);
assign g12493 = ((~g8632));
assign g17394 = ((~g16197));
assign II24494 = ((~g6301))|((~II24493));
assign g19786 = (g2040&g18879);
assign g29263 = (g28867&g8974);
assign g11624 = ((~g9062)&(~g9075)&(~g9091));
assign II15577 = ((~g7265));
assign g4532 = ((~g1515));
assign g7833 = ((~g1196));
assign g29608 = ((~g13892)&(~g29251));
assign g26597 = ((~g25443));
assign g13041 = ((~g9822))|((~g7358));
assign g11690 = ((~g9119)&(~g9124)&(~g9127));
assign g29368 = ((~g28916));
assign g17741 = ((~g13895));
assign g23381 = ((~g22013))|((~g22001));
assign g19890 = ((~II26334));
assign g13299 = ((~g8946)&(~g8979)&(~g9004));
assign g28271 = ((~II37062));
assign g8242 = ((~g2561));
assign g26954 = ((~g26549));
assign g13300 = ((~II20365));
assign g20621 = ((~II27188));
assign g17449 = (g4121&g15112);
assign g5044 = ((~g1135));
assign II28754 = ((~g21893))|((~II28753));
assign II24753 = ((~g14609))|((~II24751));
assign g23388 = ((~g21971))|((~g22336));
assign g15836 = ((~g12657))|((~g6574));
assign II13182 = ((~g995));
assign g28214 = ((~II36891));
assign g4085 = ((~g2248));
assign g20561 = ((~II27008));
assign g14471 = ((~g12155));
assign g6438 = ((~g2766));
assign II30878 = ((~g22113));
assign II20458 = ((~g10972));
assign g8579 = ((~II15787));
assign II25612 = ((~g17197));
assign g28442 = (g26114&g28163);
assign g13010 = (g8255&g10419);
assign II37868 = ((~g28321));
assign II31162 = ((~g22193));
assign g21921 = ((~g20002));
assign g20268 = (g13805&g13840&II26682);
assign g23200 = ((~II30053));
assign II40429 = ((~g30580));
assign g30879 = ((~II40889));
assign g17234 = ((~g16028)&(~g16045));
assign g4857 = ((~g2238));
assign g23682 = ((~II30838));
assign II29203 = ((~g20717));
assign g23427 = ((~g22699)&(~g21589));
assign g12052 = ((~g11379));
assign II38594 = ((~g28990));
assign II15493 = ((~g3252));
assign g24468 = ((~g24014))|((~g3806));
assign g10479 = (g7426&g5021);
assign g16935 = ((~II22885))|((~II22886));
assign g7420 = ((~g2539));
assign g19515 = ((~g18325));
assign g12152 = ((~g10378)&(~g10442)&(~g10506));
assign II34230 = ((~g25249));
assign g27054 = (g22083&g26620);
assign II23076 = ((~g13856))|((~II23074));
assign g13675 = (g7561&g12532);
assign II24545 = ((~g14263))|((~II24544));
assign g19016 = ((~II25111));
assign g23180 = ((~II29993));
assign g30857 = ((~II40823));
assign II31451 = ((~g23682));
assign II23893 = ((~g14177))|((~g9174));
assign II18632 = ((~g8850));
assign g29914 = ((~g24695)&(~g29724));
assign g24736 = ((~g23939)&(~g22830));
assign g11373 = ((~II18329));
assign II18611 = ((~g10909));
assign g28892 = (g14001&g28640);
assign g11866 = ((~g11092));
assign g17383 = ((~g16184)&(~g16238));
assign g30021 = ((~g29541)&(~g29954));
assign g16778 = ((~g15003)&(~g15161));
assign g29727 = ((~g29583)&(~g1912));
assign II15918 = ((~g6643));
assign g30841 = ((~II40775));
assign g29274 = ((~g28775));
assign g24874 = (g24060&g18899);
assign g7583 = ((~g2892));
assign g21169 = ((~g20057)&(~g20019));
assign g13370 = ((~II20466))|((~II20467));
assign g18490 = ((~g13565));
assign g22343 = ((~g20810));
assign g20842 = ((~g19441));
assign II32164 = ((~g24228));
assign g10809 = ((~g5701));
assign II40730 = ((~g30658));
assign II25044 = ((~g14273));
assign II36536 = ((~g27278));
assign g26988 = ((~g24893)&(~g26023));
assign II17030 = ((~g7053));
assign gbuf175 = (g2525);
assign II24078 = ((~g9277))|((~II24076));
assign g29154 = ((~II38205));
assign g24455 = ((~g23748))|((~g3618));
assign II23046 = ((~g9248))|((~II23045));
assign g22776 = ((~II29542));
assign g25047 = ((~g23748))|((~g7015));
assign II29918 = ((~g23068));
assign g26214 = ((~II34140));
assign g17950 = (g4979&g15574);
assign II29963 = ((~g22639));
assign g18960 = ((~II25004));
assign II28503 = ((~g21528));
assign g30081 = (g29823&g11022);
assign g22745 = (g14322&g21606);
assign II21897 = ((~g13122));
assign g25362 = (g24683&g18217);
assign g26778 = (g24929&g26516&g13626);
assign II13218 = ((~g2010));
assign g9781 = (g6369&g4044);
assign g13677 = ((~g12447));
assign g17541 = (g6298&g15222);
assign g16355 = ((~II22414));
assign g27264 = ((~g26984)&(~g26278));
assign g23713 = ((~II30881));
assign g16233 = ((~g12981))|((~g2707));
assign g10711 = (g7595&g7600&II17599);
assign II18013 = ((~g5594));
assign II22912 = ((~g15151));
assign II14550 = ((~g458));
assign g8785 = ((~II15983));
assign II21992 = ((~g13139));
assign g12914 = ((~g8952));
assign g20058 = ((~II26494));
assign g28385 = (g2124&g28041);
assign g16964 = (g7520&g15170);
assign g12221 = ((~g8421));
assign g5878 = ((~g2300));
assign g12997 = ((~g9041));
assign II37092 = ((~g28115));
assign g30002 = (g29905&g8455);
assign g12326 = ((~g10630)&(~g10663)&(~g10682));
assign II38453 = ((~g28746));
assign g18875 = ((~g15415));
assign g4570 = ((~g2253));
assign g20049 = (g17878&g3155);
assign g23030 = ((~g16970)&(~g21091));
assign II20634 = ((~g11636));
assign g28107 = ((~II36752));
assign g3981 = ((~g2217));
assign II36741 = ((~g27332));
assign g29111 = ((~g28658)&(~g17065));
assign g30807 = ((~II40673));
assign g12814 = ((~g8387)&(~g8432)&(~g8463));
assign g25217 = ((~g24758)&(~g23567));
assign g11255 = ((~II18181));
assign II20863 = ((~g12467));
assign II31625 = ((~g23661));
assign II25800 = ((~g83))|((~g18265));
assign g22107 = ((~II28649));
assign g24843 = (g21825&g23918);
assign g10302 = (g6751&g1273);
assign g8760 = (g7053&g7845);
assign g30353 = ((~II39878));
assign g20877 = ((~g3919)&(~g19830));
assign II37584 = ((~g28526));
assign g5929 = ((~g776));
assign g5759 = ((~g508));
assign g21667 = ((~g20481)&(~g6777));
assign g5740 = (g1706&g1745);
assign II40775 = ((~g30807));
assign g15812 = ((~g12711))|((~g7085));
assign g12091 = ((~II19271));
assign g20315 = ((~g17315));
assign g8417 = (g6838&g2288);
assign g25348 = (g24664&g18101);
assign g8688 = (g6945&g7858);
assign g27129 = ((~g26607)&(~g17065));
assign g22306 = ((~g20769));
assign g28239 = ((~II36966));
assign g30277 = ((~g16418)&(~g30111));
assign g15338 = (g4651&g13199);
assign g13622 = ((~II20848));
assign g19062 = ((~II25249));
assign II27972 = ((~g19163));
assign II35886 = ((~g26944));
assign g27234 = ((~II35539));
assign g25877 = ((~II33723));
assign II39038 = ((~g29551));
assign g30572 = ((~g30399));
assign g5095 = ((~g2100));
assign g23314 = ((~II30395));
assign II39997 = ((~g30248));
assign g16313 = ((~g13076));
assign II36253 = ((~g27674));
assign g24925 = (g23772)|(g23141);
assign II23625 = ((~g15898));
assign g14606 = ((~g12270));
assign g10291 = (g3366&g4620);
assign g18623 = ((~g15902)&(~g2814));
assign g27671 = (g26885&g22212);
assign g11588 = ((~II18740));
assign g13880 = (g1234&g12790);
assign g10821 = ((~II17666));
assign g11210 = ((~II18136));
assign g20323 = ((~g17330));
assign II40751 = ((~g30665));
assign g17192 = ((~II23265))|((~II23266));
assign g23190 = ((~II30023));
assign g29191 = ((~II38278));
assign II32357 = ((~g24003))|((~II32355));
assign g10288 = (g3366&g4611);
assign g17059 = ((~g15933)&(~g15913)&(~g15890));
assign g12477 = (g7822&g9128);
assign g10689 = (g3806&g5338);
assign g20062 = (g18225&g18141&II26500);
assign g27493 = ((~II35841));
assign g29236 = (g9471&g28810);
assign g6636 = ((~g1491));
assign g19172 = ((~g17635)&(~g15388));
assign g20015 = (g18183)|(g18079)|(II26455);
assign II23513 = ((~g15850));
assign g14565 = ((~g12224));
assign g25109 = ((~II32835));
assign II30113 = ((~g22790));
assign II31859 = ((~g23677));
assign g17229 = ((~g16019)&(~g16032));
assign g17097 = (g7622&g15622);
assign II38515 = ((~g28782));
assign g25187 = (g24633&g16608);
assign g12939 = ((~g8501)&(~g8516)&(~g8531));
assign II20703 = ((~g12123));
assign g24347 = ((~II31715));
assign II40313 = ((~g30505));
assign g10663 = (g7265&g5309);
assign g11794 = ((~g10974));
assign g12069 = (g7964&g8763);
assign g29139 = ((~II38160));
assign g18946 = ((~g15672));
assign g22736 = ((~II29448));
assign g23892 = ((~g23042)&(~g18604)&(~g4809));
assign g29788 = ((~g29488)&(~g29241));
assign g14249 = ((~g12034));
assign g4573 = ((~g2489));
assign gbuf7 = (g2821);
assign g25314 = ((~g24897));
assign g26689 = ((~II34674));
assign II17061 = ((~g6309))|((~II17059));
assign g18953 = ((~g15701));
assign g15783 = ((~g11643))|((~g12392));
assign g30517 = ((~II40131));
assign g13156 = ((~g8296))|((~g3618));
assign g13378 = ((~g9026)&(~g9047)&(~g9061));
assign g16866 = ((~g15840)&(~g13042));
assign II21796 = ((~g11708));
assign g22661 = ((~g21130));
assign g20977 = ((~g19784)&(~g17773));
assign II29990 = ((~g22728));
assign g8082 = ((~II15345));
assign II20359 = ((~g10838));
assign g9822 = (g7802&g6166&g1918);
assign g16468 = ((~II22506));
assign II28357 = ((~g20497));
assign g5697 = ((~g2147));
assign II34388 = ((~g25200));
assign II35834 = ((~g26792));
assign g11678 = ((~g9110)&(~g9116)&(~g9121));
assign II26285 = (g18281&g18436&g18091);
assign g11392 = ((~II18350));
assign g18833 = ((~g15237));
assign g11929 = ((~g11199));
assign g10928 = ((~g5951));
assign g20557 = ((~II26996));
assign g29425 = ((~II38656));
assign II25423 = ((~g18852));
assign g19278 = (g17998)|(g18096);
assign g27631 = ((~g26833)&(~g26053));
assign g24888 = (g24073&g18922);
assign g4107 = ((~g177));
assign g11277 = ((~II18223));
assign II20652 = ((~g12445));
assign g13200 = ((~g9592));
assign II25644 = ((~g749))|((~II25643));
assign g8378 = ((~II15580));
assign g21988 = ((~g21262)&(~g21276));
assign g22210 = ((~g21610)&(~g19932));
assign g29491 = ((~g29350));
assign g4118 = ((~g703));
assign g13079 = ((~g10855));
assign g13322 = (g5694&g11240);
assign II20813 = ((~g13265));
assign g7891 = ((~g2010));
assign g26887 = ((~g26498)&(~g5732));
assign g30643 = ((~g16200)&(~g30441));
assign II31685 = ((~g23626));
assign g30129 = (g30071&g20725);
assign g20437 = ((~g17707));
assign g25333 = ((~g24937));
assign g14171 = ((~g11979));
assign g8071 = ((~g1173));
assign g18920 = ((~g15566));
assign g21651 = ((~II28178));
assign II18653 = ((~g8971));
assign II13928 = ((~g388));
assign II14654 = ((~g3220));
assign g25488 = ((~II33316));
assign g8842 = (g6512&g5508);
assign g19159 = ((~II25358));
assign g7806 = ((~g2397));
assign II35708 = ((~g26974));
assign g29455 = ((~II38746));
assign II37632 = ((~g28372));
assign g27045 = (g23372&g26611);
assign II23445 = ((~g15808));
assign g24819 = ((~g16262)&(~g24236));
assign g26004 = ((~II33864));
assign g23084 = (g21815)|(g21810)|(g21849);
assign g5922 = ((~II14378));
assign g21001 = ((~g19818)&(~g17855));
assign gbuf41 = (g365);
assign g20717 = ((~g19165)&(~g10133));
assign g17001 = (g3254&g10694&g14144);
assign g8990 = ((~II16306));
assign II17125 = ((~g7053));
assign g25369 = ((~II33205));
assign g20146 = (g16201&g13714&g13756&II26590);
assign II29653 = ((~g21746));
assign g24957 = ((~II32719));
assign II40883 = ((~g30824));
assign II31124 = ((~g22182));
assign g8021 = ((~II15313));
assign II33479 = ((~g25032));
assign g23792 = ((~II31008));
assign g23199 = ((~II30050));
assign g26106 = ((~g23644))|((~g25354));
assign g25886 = ((~II33732));
assign g20605 = ((~II27140));
assign g23344 = ((~g23113))|((~g23099));
assign II26198 = ((~g16854));
assign g27325 = ((~g27073)&(~g26426));
assign g6205 = ((~g1243));
assign g27541 = (g24004&g27159);
assign g25145 = ((~II32913));
assign g27513 = ((~g24969)&(~g24653)&(~g26778));
assign g8215 = ((~g839));
assign g18763 = ((~g13671)&(~g11838));
assign II40661 = ((~g30635));
assign II25334 = ((~g17645));
assign g9506 = ((~g6444));
assign g16300 = (g5861&g11942);
assign g19271 = ((~II25561))|((~II25562));
assign g24800 = ((~g16211)&(~g24229));
assign II17106 = ((~g6945));
assign g18836 = ((~g13789)&(~g11967));
assign g18598 = ((~g14371)&(~g16120));
assign g15793 = (g5361&g13347);
assign g11919 = ((~g11179));
assign g26135 = ((~II34029));
assign g27098 = (g22021&g26651);
assign II24725 = ((~g6222))|((~g14626));
assign g17399 = ((~II23487));
assign g19852 = (g2052&g18920);
assign g11503 = ((~II18485));
assign g29457 = ((~II38752));
assign g30225 = (g30044&g9035);
assign g19594 = (g16935&g12555);
assign g23189 = ((~II30020));
assign g26530 = ((~g25967)&(~g17031));
assign gbuf19 = (g2858);
assign g17825 = ((~g13927));
assign g7195 = ((~II14928));
assign g8317 = ((~g3919));
assign II21868 = ((~g13134));
assign g12062 = ((~g10258)&(~g10326)&(~g10403));
assign g28690 = ((~II37617));
assign g29545 = (g29216&g29381);
assign II28235 = ((~g20153));
assign g19256 = (g17019)|(g16996)|(II25521);
assign II14502 = ((~g471));
assign g25008 = ((~g23644))|((~g5438));
assign II40086 = ((~g30265));
assign g28785 = ((~II37746));
assign g22208 = (g21654&g21057);
assign g10449 = (g3522&g4939);
assign g29064 = ((~g28327)&(~g28330));
assign II35512 = ((~g26843));
assign g28814 = ((~II37775));
assign II24399 = ((~g13936))|((~g9264));
assign g17959 = ((~II23996));
assign g21403 = (g15022&g20399);
assign g5659 = ((~g1453));
assign g27551 = ((~g4632)&(~g26882));
assign II24196 = ((~g15188))|((~II24194));
assign g20061 = (g17942)|(g18556)|(II26497);
assign g21788 = (g20117)|(g20094)|(II28305);
assign g6232 = ((~II14715));
assign II15677 = ((~g3722));
assign g26981 = (g23325&g26555);
assign g22215 = (g21285&g16940);
assign gbuf54 = (g523);
assign g29128 = ((~g28380)&(~g27783));
assign g26625 = ((~g25729));
assign g10442 = (g6945&g4922);
assign g16254 = ((~g13060));
assign II31556 = ((~g23439));
assign g14497 = ((~g12994));
assign g15453 = (g6898&g12811);
assign g26458 = ((~g25343))|((~g65));
assign g18297 = ((~g14292));
assign g30587 = ((~II40313));
assign g28788 = ((~g28476)&(~g27984));
assign II33352 = ((~g24443));
assign g4578 = ((~g2772));
assign II14343 = ((~g3219));
assign g28609 = ((~g27839));
assign g5852 = ((~g121));
assign g16239 = (g5700&g11887);
assign g25972 = (g24859&g12042);
assign g19106 = (g14863&g18735&g18765&g16395);
assign II24187 = ((~g6177))|((~II24186));
assign g29953 = (g29791&g28967);
assign g24416 = ((~II31922));
assign g20399 = ((~g17563));
assign g30108 = (g29877&g11401);
assign II18641 = ((~g8871));
assign g11581 = ((~II18719));
assign g28016 = ((~II36521));
assign g8076 = ((~g1524));
assign g13755 = (g7347&g12551);
assign g21808 = (g18688)|(g20282)|(g20271)|(g18650);
assign g11510 = ((~II18506));
assign II25561 = ((~g56))|((~II25560));
assign gbuf206 = (g2640);
assign g19950 = ((~g18598));
assign g30923 = (g30789&g22338);
assign g10589 = (g3774&g5201);
assign g9887 = (g6232&g4095);
assign g19147 = ((~II25338));
assign g23482 = ((~g22197));
assign g28883 = ((~II37854));
assign g28323 = (g8580&g27838);
assign g19701 = (g4234&g17511);
assign g30040 = ((~g29914));
assign g15822 = ((~g12611))|((~g6369));
assign II33810 = ((~g25646));
assign g8543 = (g3722&g2330);
assign II24340 = ((~g14438))|((~II24338));
assign g27144 = ((~g23451)&(~g26052));
assign g21198 = (g19534&g14601);
assign g28726 = (g28578&g16767);
assign g25386 = ((~II33219));
assign g20283 = (g18708&g14991&g16395);
assign g16459 = (g5997&g12174);
assign g18302 = ((~II24307))|((~II24308));
assign II30320 = ((~g22773));
assign g23573 = (g3937&g22451);
assign II13980 = ((~g2448));
assign II32460 = ((~g18247))|((~g24057));
assign g21855 = ((~g17919))|((~g19188))|((~g19193));
assign g27384 = ((~g27140));
assign g13502 = (g6036&g12264);
assign g29985 = (g29897&g8363);
assign g14290 = ((~g12049));
assign g3996 = ((~g3073));
assign g18881 = ((~g15446));
assign g7706 = ((~g1004));
assign II40578 = ((~g30702));
assign g28733 = ((~g28424)&(~g27909));
assign g29446 = ((~II38719));
assign g29254 = ((~II38363));
assign g17172 = (g7730&g14230);
assign g10500 = ((~g7962));
assign g7730 = ((~g2478));
assign g22234 = ((~g21670)&(~g19976));
assign g4879 = ((~g2803));
assign II31691 = ((~g24053));
assign g29569 = ((~g28708)&(~g29174));
assign gbuf162 = (g1915);
assign g23637 = (g4194&g22540);
assign g6081 = ((~II14590));
assign g19357 = ((~II25762))|((~II25763));
assign g29441 = ((~II38704));
assign g13536 = ((~g12711))|((~g3722));
assign g20303 = ((~g17285));
assign II24640 = ((~g14390))|((~II24639));
assign II15565 = ((~g6838));
assign II36479 = ((~g27504));
assign g5866 = ((~g1426));
assign g4655 = ((~g1273));
assign II16027 = ((~g3806));
assign g20374 = ((~g17482));
assign g23017 = ((~g21696))|((~g2052));
assign II29948 = ((~g22549));
assign II13161 = ((~g308));
assign g27036 = ((~g26070));
assign g27240 = (g26905&g22241);
assign II20517 = ((~g12425));
assign g27938 = (g14053&g27443);
assign II24318 = ((~g6832))|((~II24317));
assign g19719 = (g4298&g17548);
assign g29869 = ((~g29679));
assign g10156 = (g7015&g1801);
assign g27197 = ((~II35428));
assign g20624 = ((~II27197));
assign g12433 = ((~g2879))|((~g10778));
assign g9746 = (g7085&g3984);
assign II28115 = ((~g20493));
assign II38450 = ((~g28745));
assign g26090 = ((~g25518)&(~g25560));
assign g21517 = (g9711&g20461);
assign II17043 = (g5886&g6040&g5199&g5200);
assign g8177 = ((~g3043));
assign g8748 = ((~II15938));
assign II29712 = ((~g21786));
assign g22259 = ((~II28833));
assign II37986 = ((~g28529));
assign g11803 = ((~g10994));
assign g10354 = ((~g7815))|((~g3834));
assign g9371 = ((~II16581));
assign g5700 = ((~g3088));
assign g18604 = ((~g13582));
assign g21654 = (g14053&g14502&g19907&II28181);
assign g28458 = ((~II37415));
assign g23266 = ((~II30251));
assign g22530 = ((~II29080));
assign g21514 = ((~II28047));
assign g13635 = ((~II20863));
assign g27572 = ((~g26911)&(~g24717));
assign g5830 = ((~II14280));
assign II18761 = ((~g9005));
assign g15829 = (g7857&g13400);
assign II22651 = ((~g14677));
assign g5081 = ((~g1960));
assign g24440 = (g24168&g13649);
assign g16712 = ((~g14863));
assign g22563 = ((~II29125));
assign g27079 = (g5044&g26401);
assign g19565 = (g8126&g17275);
assign g11932 = ((~g11209));
assign g20089 = (g17969&g9160);
assign g20288 = ((~g17255));
assign II32193 = ((~g23513));
assign g15994 = ((~g12555));
assign g4504 = ((~g850));
assign g5437 = ((~II13999));
assign g8194 = ((~g152));
assign g9939 = (g7230&g4176);
assign g26031 = ((~g25273)&(~g22777));
assign g11799 = ((~g9520)&(~g9631)&(~g9759));
assign II35446 = ((~g26762));
assign g10065 = (g5512&g1798);
assign g9006 = ((~II16328));
assign g15950 = ((~g12711))|((~g7085));
assign II18584 = ((~g8677));
assign g29947 = (g29785&g28911);
assign g8627 = ((~II15815));
assign g24498 = ((~g15324)&(~g23777));
assign g16336 = (g5662&g13300);
assign II15946 = ((~g5692));
assign II36876 = ((~g27986));
assign II39243 = ((~g29694));
assign g24095 = ((~g22362));
assign g20330 = ((~g17354));
assign g28967 = ((~II37934));
assign g25327 = ((~II33157));
assign g10458 = (g7195&g1970);
assign g30885 = ((~II40907));
assign II29049 = ((~g21750));
assign g24175 = ((~g22592));
assign g21329 = (g9161&g20328);
assign g10534 = (g7391&g2664);
assign II20694 = ((~g13346));
assign g21380 = (g15096&g20380);
assign g3337 = ((~g309));
assign g14609 = ((~g12271));
assign g24271 = ((~II31487));
assign g21494 = (g6632&g19792);
assign g22428 = ((~II28972));
assign II30614 = ((~g22031));
assign II39818 = ((~g30215));
assign g13000 = (g7973&g10357);
assign g23944 = (g7570&g23103);
assign II17370 = ((~g3900));
assign II21723 = ((~g13088));
assign g25192 = (g24711&g20790);
assign g24380 = ((~II31814));
assign g21011 = ((~g19841)&(~g17902));
assign g18314 = ((~g14322));
assign II27257 = ((~g19431));
assign g20080 = (g18586&g18537&II26508);
assign g27942 = ((~II36407));
assign II18103 = ((~g7391));
assign II34650 = ((~g26172));
assign g28097 = ((~II36724));
assign g15699 = (g5278&g13283);
assign II23836 = ((~g13559));
assign g5072 = ((~g1757));
assign g20486 = (g17281&g11859);
assign g22054 = ((~g21319)&(~g19586));
assign II32402 = ((~g24036))|((~II32400));
assign g23286 = ((~II30311));
assign g27594 = ((~g27175)&(~g17001));
assign g22163 = ((~g21439)&(~g19771));
assign g15803 = ((~g13375))|((~g12354));
assign g11825 = ((~g11025));
assign II30797 = ((~g22087));
assign g25156 = ((~II32946));
assign g12212 = ((~g8408));
assign II32597 = ((~g23938))|((~II32595));
assign II28726 = ((~g21887))|((~g13519));
assign g24327 = ((~II31655));
assign g19035 = ((~II25168));
assign g24470 = ((~g23984))|((~g3650));
assign g19171 = ((~g17616)&(~g15356));
assign g17446 = (g6284&g16011);
assign g16907 = (g7335&g15017);
assign g30894 = ((~II40934));
assign g5382 = ((~g2117));
assign g30951 = (g30934&g20833);
assign g14773 = (g7915&g13141);
assign g26692 = ((~II34683));
assign g24114 = ((~g22451));
assign g20456 = ((~g17799));
assign II32669 = ((~g18247))|((~II32668));
assign g14039 = (g7688&g12931);
assign g18986 = ((~II25050));
assign g28306 = ((~II37167));
assign II17685 = ((~g6630));
assign g21396 = (g9407&g20392);
assign g5887 = ((~g2581));
assign g29420 = ((~II38641));
assign g25320 = ((~g21219))|((~g14529))|((~g10714))|((~g24595));
assign II37059 = ((~g28099));
assign g17471 = ((~II23559));
assign II16065 = ((~g7936));
assign g12972 = ((~g9013));
assign II18542 = ((~g10968));
assign g8569 = ((~II15771));
assign g11264 = ((~II18205))|((~II18206));
assign g21158 = (g19505&g14459);
assign g23285 = ((~II30308));
assign II29603 = ((~g21051));
assign g4079 = ((~g2227));
assign g27988 = ((~II36465));
assign g23617 = (g22810&g20382);
assign g24278 = ((~II31508));
assign II26966 = ((~g17051));
assign g6039 = ((~g2348));
assign II38321 = ((~g29113));
assign g11638 = ((~II18824));
assign II35883 = ((~g26781));
assign g9064 = (g6713&g7632);
assign g12537 = ((~g8681));
assign g29331 = ((~II38510));
assign II14973 = ((~g2006));
assign g21594 = ((~II28123));
assign g14252 = ((~g12035));
assign g26793 = ((~II34916));
assign g29993 = (g29897&g8411);
assign g10612 = (g3494&g5238);
assign II33246 = ((~g24890));
assign g20538 = (g18656&g14837&g13657&g16189);
assign g21627 = ((~g19330));
assign II20493 = ((~g10934));
assign g16595 = (g15942)|(g14725);
assign g27027 = (g21991&g26598);
assign g11742 = ((~g10883));
assign g11098 = ((~II18010));
assign II35036 = ((~g26154))|((~II35034));
assign II39339 = ((~g29748))|((~g29741));
assign g23827 = ((~II31053));
assign II14857 = ((~g626));
assign g16113 = ((~g11903));
assign II13953 = ((~g1075));
assign g24479 = ((~g23593)&(~g22516));
assign g29758 = ((~g16335)&(~g29619));
assign g22790 = ((~II29556));
assign II28061 = ((~g19178));
assign g13110 = (g10693&g2883&g7562&g10711);
assign II18265 = ((~g3722));
assign g27020 = (g22069&g26588);
assign g30952 = ((~II41065))|((~II41066));
assign II38626 = ((~g29297));
assign g3941 = ((~g455));
assign II32889 = ((~g24568));
assign g26605 = ((~g25661));
assign g27969 = ((~g27361));
assign II18241 = ((~g6713));
assign g22728 = ((~II29426));
assign g5796 = ((~II14238));
assign g29657 = ((~II39089));
assign g20442 = ((~g17738));
assign g22490 = ((~II29036));
assign g22881 = ((~g8287))|((~g21689));
assign g26261 = (g25895&g9443);
assign II21933 = ((~g11723));
assign II32140 = ((~g24216));
assign g12859 = ((~g8901));
assign II27083 = ((~g19208));
assign g13922 = ((~g11831));
assign II39916 = ((~g30293));
assign II21274 = ((~g11653));
assign g13856 = ((~g11759));
assign g25515 = ((~II33343));
assign g16003 = (g12013&g10826);
assign g17563 = ((~II23651));
assign g17530 = (g4263&g15207);
assign g8203 = ((~g173));
assign g26548 = ((~II34505));
assign g28250 = ((~II36999));
assign g22620 = ((~II29206));
assign g30774 = ((~II40584));
assign II34032 = ((~g25520));
assign g29775 = ((~g29476)&(~g29217));
assign g25177 = ((~II33009));
assign g4082 = ((~g2246));
assign g9116 = (g7265&g7745);
assign II19507 = ((~g10606));
assign g7541 = ((~g2180));
assign g29373 = ((~g28945));
assign g19468 = ((~g17216));
assign II20032 = ((~g10003))|((~II20031));
assign g23630 = (g4165&g22527);
assign g18619 = ((~II24732));
assign g26291 = (g25899&g9524);
assign g21687 = (g3398&g20516);
assign g6675 = ((~g458));
assign g27249 = (g27065&g16775);
assign g5508 = ((~II14014));
assign g26471 = ((~II34433));
assign g27225 = ((~II35512));
assign g23291 = ((~II30326));
assign g19450 = (g14837)|(g16682);
assign g26906 = ((~g25772))|((~g26327))|((~g25648))|((~g25708));
assign g16344 = (g5896&g11970);
assign g24809 = (g15694&g24159);
assign II19500 = ((~g10424));
assign g22556 = (g20904&g17523);
assign g3247 = ((~II13137));
assign g25141 = ((~II32901));
assign g23087 = ((~g21651));
assign g13394 = ((~II20493));
assign g11179 = ((~II18097));
assign g23230 = ((~II30143));
assign g9819 = ((~II16857));
assign II25783 = ((~g18207))|((~II25781));
assign g15859 = ((~g13378));
assign g8484 = (g6232&g186);
assign gbuf215 = (g2594);
assign g29770 = ((~g29471)&(~g29196));
assign II18025 = ((~g6574));
assign g13207 = ((~g9666));
assign II14424 = ((~g117));
assign g10431 = (g6643&g4891);
assign g20397 = ((~g17557));
assign II23878 = ((~g14001))|((~g9187));
assign g25281 = (g5606&g24815);
assign g10541 = (g7426&g5138);
assign g12251 = ((~g8440));
assign g12498 = ((~g8637));
assign g27912 = ((~II36371));
assign II17709 = ((~g6894));
assign g13247 = (g298&g11032);
assign gbuf39 = (g352);
assign g17579 = ((~II23667));
assign g12825 = ((~II19886));
assign II29456 = ((~g20999));
assign g15739 = (g5318&g13303);
assign II37277 = ((~g28146));
assign g26789 = ((~g26046)&(~g10238));
assign g14024 = ((~II21045));
assign II23992 = ((~g13564));
assign II31253 = ((~g22231));
assign g27716 = ((~II36159));
assign II26348 = (g18448&g14028&g14102);
assign g4351 = ((~g709));
assign g18866 = ((~g13834)&(~g12069));
assign g24143 = ((~g22503));
assign g29808 = ((~II39276));
assign g28838 = (g5866&g28496);
assign II22542 = ((~g14954));
assign g24389 = ((~II31841));
assign g20898 = ((~g19636)&(~g17464));
assign g21196 = (g19329&g19313&II27761);
assign g8512 = (g7085&g2318);
assign g7691 = ((~g1696));
assign II40149 = ((~g30358));
assign g23461 = ((~g22841)&(~g21707));
assign II27140 = ((~g19690));
assign II25763 = ((~g17882))|((~II25761));
assign g30465 = (g30175&g11252);
assign II35376 = ((~g26336));
assign g11592 = ((~II18752));
assign g28046 = ((~II36592))|((~II36593));
assign g30276 = ((~g16415)&(~g30110));
assign g4315 = ((~g2773));
assign g9816 = ((~II16854));
assign II38881 = ((~g29187));
assign g23544 = (g5992&g22868);
assign II26934 = ((~g17341));
assign g27959 = ((~II36426));
assign g23360 = ((~g21980))|((~g21975));
assign II29183 = ((~g21792));
assign II34029 = ((~g25520));
assign g24789 = (g9711&g24141);
assign g18011 = (g5058&g15606);
assign g17275 = ((~II23361));
assign g30785 = ((~g30618)&(~g22387));
assign g26724 = ((~II34779));
assign g30818 = ((~II40706));
assign g4734 = ((~g11));
assign g16023 = ((~g12699));
assign II39340 = ((~g29748))|((~II39339));
assign g18395 = ((~II24416))|((~II24417));
assign II31088 = ((~g22172));
assign g5663 = ((~g3179));
assign g12445 = ((~II19611));
assign g29147 = ((~II38184));
assign g21143 = (g19494&g18121&g14309);
assign g26516 = ((~g25320));
assign g28433 = (g28133&g9212);
assign g13327 = ((~II20398));
assign g10875 = ((~II17734));
assign g22361 = ((~g20246)&(~g21822));
assign g29849 = ((~g29671));
assign II13925 = ((~g376));
assign g29547 = (g29219&g29382);
assign g27496 = ((~g27185)&(~g25178));
assign II23430 = ((~g13494));
assign g25711 = ((~II33539));
assign II39414 = ((~g29658));
assign g24768 = (g9569&g24122);
assign g24526 = ((~g23848)&(~g22719));
assign II24006 = ((~g7548))|((~II24005));
assign II34997 = ((~g26482));
assign g15109 = ((~II21429));
assign g8264 = ((~II15460));
assign II36296 = ((~g27626));
assign g29381 = ((~g28983));
assign g19752 = (g2013&g18859);
assign II38003 = ((~g28529));
assign II27170 = ((~g20396));
assign II27308 = ((~g19401));
assign II16092 = ((~g5402));
assign g18842 = ((~g15268));
assign g21260 = (g19608&g14976);
assign II20574 = ((~g12534));
assign g26972 = (g14033&g26223);
assign g19553 = (g7990&g17237);
assign g23721 = (g4430&g22600);
assign g26315 = ((~II34277));
assign g27682 = ((~g26801)&(~g10238));
assign II38181 = ((~g28899));
assign g17422 = ((~II23510));
assign g27102 = ((~II35283));
assign II29872 = ((~g21364));
assign g8015 = ((~g2941));
assign g10691 = (g7391&g2691);
assign II29246 = ((~g20922));
assign g19772 = (g4504&g17661);
assign g23125 = ((~II29872));
assign g11997 = ((~g11309));
assign g23508 = ((~II30552));
assign g24865 = ((~II32535));
assign g8433 = (g6232&g249);
assign g25203 = ((~g24978))|((~g3462));
assign g4275 = ((~g1556));
assign II30766 = ((~g22077));
assign g21138 = (g19484&g14347);
assign gbuf113 = (g1221);
assign g18794 = ((~g13701)&(~g11880));
assign II37110 = ((~g28067));
assign g6018 = ((~g894));
assign g20951 = ((~g19743)&(~g17675));
assign g22335 = ((~g20802));
assign g13614 = ((~g11690));
assign g10898 = ((~II17771));
assign g25026 = ((~g23803))|((~g7265));
assign g24501 = ((~g15339)&(~g23790));
assign g10973 = ((~II17872));
assign g23766 = ((~II30962));
assign g13788 = (g6897&g12553);
assign g8949 = ((~II16255));
assign II37119 = ((~g28089));
assign g21290 = (g9356&g20278);
assign g11728 = ((~g9968))|((~g3834));
assign g6139 = ((~II14654));
assign g29170 = ((~g28844)&(~g28399));
assign g5415 = ((~II13959));
assign g19523 = ((~g16814));
assign g20298 = ((~g17278));
assign g26404 = (g5047&g25714);
assign II32308 = ((~g17903))|((~g23973));
assign II17884 = ((~g8031));
assign g28772 = ((~g28454)&(~g27949));
assign II40542 = ((~g30695));
assign g21120 = (g19484)|(g16515)|(g14071);
assign g23149 = ((~II29900));
assign g27307 = ((~g27047)&(~g26386));
assign gbuf158 = (g1948);
assign g18639 = ((~g14570)&(~g16230));
assign g21470 = ((~g20512)&(~g16417));
assign II40521 = ((~g30689));
assign g9641 = ((~II16744));
assign g24508 = ((~g15392)&(~g23825));
assign g13436 = ((~II20607));
assign g30811 = ((~II40685));
assign II32626 = ((~g23969))|((~II32624));
assign g12114 = ((~g10324)&(~g10402)&(~g10466));
assign g13547 = ((~g12565))|((~g3254));
assign g5399 = ((~II13913));
assign g5771 = ((~II14219));
assign g9128 = ((~II16432));
assign g26568 = ((~g25546));
assign g28986 = (g14390&g28652);
assign II25123 = ((~g18890));
assign g21078 = (g20099&g14309&g14402);
assign g24751 = (g9427&g24105);
assign g19308 = ((~II25654))|((~II25655));
assign g8483 = (g6838&g2306);
assign g15660 = ((~g13401))|((~g12354));
assign g23420 = ((~g23089));
assign g18351 = ((~g13741));
assign g27721 = (g27579&g20655);
assign g4159 = ((~g1537));
assign II37939 = ((~g28501));
assign II40555 = ((~g30699));
assign g19057 = ((~II25234));
assign g26160 = ((~g25951)&(~g16162));
assign g15254 = ((~II21537));
assign II32137 = ((~g24215));
assign g22060 = ((~g21325)&(~g19592));
assign II39386 = ((~g29710))|((~II39384));
assign g24437 = (g24153&g13637);
assign II19598 = ((~g9215));
assign g5298 = ((~g1828));
assign g27805 = ((~II36264));
assign g28347 = ((~II37238));
assign g17049 = ((~II23028))|((~II23029));
assign II35750 = ((~g26928));
assign g29217 = (g15274&g28775);
assign g25560 = (g24494&g17764);
assign II34020 = ((~g25940));
assign g16128 = ((~g12860));
assign g15317 = ((~II21586));
assign g23777 = (g22949&g9528);
assign g15899 = ((~g12657))|((~g6783));
assign g22803 = ((~II29591));
assign g22844 = ((~g21865))|((~g21860))|((~g21857));
assign g3954 = ((~g842));
assign II20407 = ((~g9027));
assign g15234 = (g4436&g13183);
assign g28928 = ((~II37897));
assign g7575 = ((~g2984)&(~g2985));
assign g10314 = (g5512&g1819);
assign II40913 = ((~g30774));
assign g19680 = ((~g16971));
assign g28411 = (g7809&g27872);
assign g30054 = ((~g29964)&(~g16336));
assign II40242 = ((~g30379));
assign g22784 = ((~g16075)&(~g20885));
assign g21962 = ((~II28512));
assign g20629 = ((~II27212));
assign g30487 = ((~g14114)&(~g30221));
assign g9099 = (g5512&g7694);
assign g5940 = ((~g1633));
assign II36126 = ((~g27553));
assign g26864 = ((~II35031));
assign II30182 = ((~g22683));
assign g23401 = ((~g22566)&(~g21452));
assign g19871 = (g14086&g18275&II26311);
assign g21816 = (g19138)|(g19681)|(g16743);
assign g9812 = ((~II16850));
assign g30837 = ((~II40763));
assign g24560 = ((~II32098));
assign g22189 = ((~g19899)&(~g21622));
assign g8513 = (g6838&g2324);
assign g16025 = ((~g12705));
assign g11542 = ((~II18602));
assign gbuf104 = (g1250);
assign II16462 = ((~g5438));
assign g11838 = (g6205&g8659);
assign g28217 = ((~II36900));
assign g8561 = (g3566&g1582);
assign g22311 = (g21782&g12346);
assign g3722 = ((~II13221));
assign g25306 = ((~II33136));
assign g8693 = ((~II15893));
assign g10744 = ((~g3710))|((~g7230));
assign II35076 = ((~g26532));
assign g23581 = ((~II30663));
assign g25236 = ((~g24792)&(~g23609));
assign g4894 = ((~g585));
assign g22711 = ((~II29389));
assign g27451 = ((~II35791));
assign g11974 = ((~g10105)&(~g10194)&(~g10279));
assign g27151 = ((~g26401));
assign g17314 = ((~g16110));
assign g22506 = ((~II29052));
assign II31874 = ((~g23720));
assign g10664 = ((~g8168));
assign g18781 = ((~g13675)&(~g11851));
assign II25162 = ((~g16863));
assign II23348 = ((~g15786));
assign g29197 = ((~g15031)&(~g28893));
assign g24334 = ((~II31676));
assign g21862 = ((~g18195))|((~g19203))|((~g19211));
assign g27203 = ((~II35446));
assign g24391 = ((~II31847));
assign g26810 = ((~g15259)&(~g26271));
assign g26233 = (g4340&g25476);
assign g26017 = ((~II33903));
assign g8851 = ((~II16095));
assign g17735 = (g4614&g15396);
assign II36362 = ((~g27667));
assign g15904 = ((~g11644));
assign g14186 = ((~g11987));
assign g5278 = ((~g2676));
assign II32860 = ((~g23803));
assign II33205 = ((~g24833));
assign g9662 = (g6369&g3954);
assign II40260 = ((~g30339));
assign g30323 = ((~II39812));
assign g20982 = ((~g19796)&(~g17796));
assign g25903 = ((~g24950));
assign II24438 = ((~g15022))|((~II24436));
assign g27727 = (g27414&g19301);
assign g5366 = ((~g2878));
assign II30371 = ((~g22749));
assign g28649 = ((~g27973));
assign g15850 = ((~g12711))|((~g6838));
assign g21949 = ((~II28473));
assign II15839 = ((~g5613));
assign g28021 = ((~II36530));
assign g29803 = ((~II39261));
assign II30065 = ((~g22621));
assign g15519 = (g4879&g12840);
assign g17341 = ((~g16138)&(~g16185));
assign g28114 = ((~II36769));
assign g29933 = ((~II39401));
assign g8867 = ((~II16123));
assign g21103 = (g20273&g12228);
assign II33145 = ((~g24997));
assign g30349 = ((~II39870));
assign g14118 = ((~g10767))|((~g12510));
assign II28047 = ((~g20481));
assign II33554 = ((~g24511));
assign g10671 = (g7391&g5315);
assign g30391 = (g30233&g8958);
assign g12084 = ((~g11425));
assign g24364 = ((~II31766));
assign g29688 = ((~g29575)&(~g29346));
assign g19911 = (g2740&g18954);
assign II30344 = ((~g22838));
assign g28653 = ((~g27999));
assign g29560 = (g29227&g29391);
assign g7862 = ((~g1859));
assign g11735 = ((~g10859));
assign II19747 = ((~g8726));
assign g6024 = ((~II14489));
assign g14831 = ((~g11828));
assign g30536 = ((~II40188));
assign g26995 = (g21991&g26563);
assign g21363 = (g15022&g20364);
assign g4175 = ((~g1836));
assign II40215 = ((~g30501));
assign g27373 = ((~II35695));
assign g27343 = ((~g27099)&(~g26477));
assign g15047 = (g4143&g13162);
assign g21572 = (g20542)|(g19505)|(g16507);
assign II39377 = ((~g15942))|((~II39375));
assign g10434 = (g6486&g605);
assign g30562 = ((~II40266));
assign g14725 = ((~II21282));
assign g5614 = ((~g1894));
assign g9968 = (g7815&g6193&g2612);
assign II18962 = ((~g9159));
assign g16463 = ((~g13004))|((~g3018));
assign g21344 = (g9150&g20345);
assign g8900 = ((~II16176));
assign II18563 = ((~g8897));
assign g5611 = ((~g1481));
assign II29274 = ((~g20934));
assign II28479 = ((~g21795));
assign g5334 = ((~II13868));
assign g23303 = ((~II30362));
assign g22359 = ((~g20819));
assign g18647 = (g14895&g16142&g16243);
assign g16222 = (g5794&g11883);
assign II29797 = ((~g21432));
assign g5634 = ((~g1895));
assign II14621 = ((~g2533));
assign g8527 = (g3722&g2321);
assign g26334 = (g4775&g25596);
assign g19854 = (g18038&g16128);
assign g25685 = ((~II33511));
assign g4870 = ((~g2778));
assign g30335 = ((~II39840));
assign g7649 = ((~g404));
assign II21289 = ((~g12434));
assign g24890 = (g23639)|(g23144);
assign II27062 = ((~g19217));
assign g24939 = ((~g23660));
assign g11493 = ((~II18455));
assign g20833 = ((~II27422));
assign g26801 = ((~g26171)&(~g25461));
assign g19239 = ((~II25492));
assign II24576 = ((~g6216))|((~II24575));
assign g18109 = ((~II24124))|((~II24125));
assign g8101 = ((~g2997));
assign g5156 = ((~g1267));
assign g4888 = ((~g578));
assign g30496 = (g30195&g11428);
assign g21320 = (g9310&g20316);
assign II19722 = ((~g10332));
assign g26622 = ((~g25714));
assign II25280 = (g18656&g18670&g18720);
assign II14442 = ((~g2165));
assign g8328 = (g6314&g225);
assign g30705 = ((~g14097)&(~g30393));
assign g12373 = ((~II19533));
assign g12646 = ((~g8788));
assign g24294 = ((~II31556));
assign g11526 = ((~II18554));
assign g28179 = ((~II36848));
assign g11036 = ((~II17951));
assign II29509 = ((~g21018));
assign II23132 = ((~g9391))|((~II23131));
assign g20217 = (g14863&g18735&g16266&g16313);
assign g11578 = ((~II18710));
assign g5631 = ((~g767));
assign II26923 = ((~g17302));
assign II30938 = ((~g22130));
assign II16993 = ((~g6643));
assign g13565 = ((~g12192));
assign II16457 = ((~g7936));
assign II14734 = ((~g135));
assign g29356 = ((~g29120));
assign II29223 = ((~g20916));
assign g8829 = ((~II16059));
assign g15064 = (g4174&g13163);
assign g25129 = ((~g23536)&(~g22383));
assign g28475 = (g28141&g9498);
assign g5315 = ((~g2660));
assign g28867 = ((~g28418));
assign g25579 = ((~II33402));
assign II27684 = ((~g20526));
assign II38275 = ((~g28987));
assign g29202 = ((~g28897)&(~g28450));
assign g27088 = (g23381&g26645);
assign II30875 = ((~g22112));
assign g25449 = ((~g24660));
assign g23848 = (g18226&g23045);
assign g13706 = ((~g12443));
assign g10514 = (g3522&g5067);
assign II13931 = ((~g1048));
assign II34683 = ((~g26364));
assign g25934 = ((~g25000))|((~g7265));
assign II23209 = ((~g13867))|((~II23207));
assign g29625 = (g29189&g11472);
assign g23643 = (g17802&g22991);
assign II26599 = (g18708&g14991&g13724);
assign II25165 = ((~g16831));
assign g27131 = ((~g26630)&(~g17100));
assign g4483 = ((~g712));
assign g29406 = ((~g28838)&(~g28387));
assign g11571 = ((~II18689));
assign g27917 = ((~g16220)&(~g27660));
assign II28159 = ((~g20067));
assign II30917 = ((~g22806));
assign g30781 = ((~II40611));
assign II21398 = ((~g13021));
assign g11915 = ((~g9940)&(~g10075)&(~g10167));
assign g11941 = ((~g11216));
assign g27984 = (g4721&g27486);
assign g9779 = (g3410&g4038);
assign II28107 = ((~g20025));
assign g30753 = ((~II40537));
assign g26529 = ((~g25962)&(~g17001));
assign g23093 = ((~g17056)&(~g21155));
assign g8181 = ((~g48));
assign g29223 = ((~g28962)&(~g28480));
assign g4591 = ((~g2870));
assign g26766 = (g14725&g26521);
assign g11780 = ((~g9440)&(~g9519)&(~g9630));
assign II23034 = ((~g9232))|((~g13864));
assign g16539 = (g15880)|(g14657);
assign g19933 = ((~g18548));
assign g29637 = ((~II39029));
assign g9890 = (g6232&g4104);
assign g5803 = ((~g117));
assign g29500 = ((~II38821))|((~II38822));
assign II30623 = ((~g22033));
assign II31565 = ((~g24001));
assign II34782 = ((~g26385));
assign g29086 = ((~II38059));
assign g3240 = ((~II13116));
assign II34425 = ((~g25270));
assign g25205 = ((~g24989))|((~g3618));
assign g8312 = ((~g3833));
assign g28465 = (g28141&g9416);
assign g4200 = ((~II13366));
assign II27318 = ((~g19457));
assign g11607 = (g5871&g8360);
assign g13183 = ((~g9416));
assign g30453 = (g30167&g11179);
assign g26026 = (g25431&g24929);
assign g23492 = ((~II30536));
assign g27622 = ((~g27174));
assign g23888 = (g18358&g23069);
assign II21747 = ((~g13116));
assign g13058 = ((~g9534))|((~g6678));
assign g23225 = ((~II30128));
assign II21426 = ((~g11661));
assign II26819 = ((~g17226));
assign II40236 = ((~g30373));
assign II24278 = ((~g6284))|((~g13918));
assign g22690 = (g21939&g12837);
assign II24158 = ((~g9407))|((~II24156));
assign g15652 = ((~II21905));
assign II23472 = ((~g13510));
assign II23084 = ((~g13879))|((~II23082));
assign II38704 = ((~g29405));
assign g28644 = ((~g27946));
assign II22945 = ((~g15188))|((~g14015));
assign g9117 = (g5556&g7748);
assign g13263 = ((~g10090));
assign g16570 = ((~g15904)&(~g15880)&(~g14630));
assign g15393 = ((~II21655));
assign g10838 = ((~II17685));
assign g30868 = ((~II40856));
assign g17294 = ((~II23380));
assign g19266 = (g17148)|(g17123)|(II25549);
assign g26664 = ((~g25346)&(~g17138));
assign g4806 = ((~g1514));
assign g19627 = (g633&g18806);
assign g12781 = ((~g8329)&(~g8386)&(~g8431));
assign g27006 = (g21991&g26579);
assign g30529 = ((~II40167));
assign g9104 = (g6713&g7709);
assign g28668 = ((~g27736)&(~g10024));
assign II14516 = ((~g3215));
assign g3617 = ((~g1686));
assign g29798 = ((~II39246));
assign g14000 = ((~g11890));
assign g7391 = ((~II14984));
assign g27864 = ((~g27632)&(~g1219));
assign g23008 = ((~g21498));
assign gbuf122 = (g1562);
assign g8594 = ((~g6623));
assign II37572 = ((~g28524));
assign g22681 = ((~g21144));
assign g22129 = ((~g21392)&(~g19704));
assign g27136 = ((~g26196));
assign g13196 = ((~g9528));
assign g7845 = ((~g1860));
assign II31727 = ((~g23602));
assign g28893 = (g28612&g9245);
assign g4026 = ((~g727));
assign gbuf129 = (g1661);
assign g19298 = (g18053)|(g18147);
assign g15682 = ((~II21933));
assign II18599 = ((~g8933));
assign g28286 = ((~II37107));
assign g25850 = ((~II33692));
assign g5426 = ((~II13990));
assign g26964 = ((~II35153));
assign g29747 = ((~g29583)&(~g1916));
assign g20418 = ((~II26843));
assign g13998 = (g7972&g12907);
assign g20367 = ((~g17454));
assign g5769 = (g1012&g1081);
assign g13405 = ((~II20514));
assign g30638 = ((~g16159)&(~g30411));
assign g18626 = ((~g16463)&(~g7549));
assign g25111 = ((~g23874));
assign g19975 = ((~g18007));
assign g17859 = ((~II23920));
assign g4452 = ((~g17));
assign g29505 = ((~II38842))|((~II38843));
assign g3304 = ((~II13161));
assign g26226 = ((~II34162));
assign g19983 = (g5352&g18432);
assign g8572 = (g3722&g2276);
assign g25890 = ((~g4985)&(~g15074)&(~g25099));
assign g5204 = ((~g2463));
assign II32325 = ((~g23982))|((~II32323));
assign g4829 = ((~g1956));
assign g7085 = ((~II14900));
assign g30138 = (g30069&g20816);
assign II34986 = ((~g26160));
assign II31071 = ((~g22168));
assign g30406 = ((~g30009)&(~g30138));
assign g26842 = (g5689&g26275);
assign g16007 = ((~g12647));
assign II16987 = ((~g6079));
assign II13116 = ((~g14));
assign g16349 = (g5902&g11984);
assign g11859 = ((~g11088));
assign g20498 = ((~II26947));
assign g30171 = ((~g30019));
assign g26897 = ((~g26513)&(~g5790));
assign g4032 = ((~g843));
assign g19826 = (g2727&g18903);
assign g24422 = ((~II31940));
assign II18784 = ((~g9067));
assign II30257 = ((~g22718));
assign II38486 = ((~g28763));
assign g22403 = ((~g21602));
assign g29385 = ((~g29005));
assign g28958 = (g14268&g28649);
assign II17159 = ((~g3900));
assign II22755 = ((~g14650));
assign II35844 = ((~g26808));
assign g7923 = ((~II15245))|((~II15246));
assign g5021 = ((~g2806));
assign II30038 = ((~g22673));
assign g17688 = ((~II23772));
assign g25016 = ((~g23748))|((~g7015));
assign g11988 = ((~g10123)&(~g10211)&(~g10298));
assign g25779 = ((~II33614));
assign II38746 = ((~g29270));
assign II26871 = ((~g17235));
assign g9921 = (g7162&g4153);
assign II17209 = ((~g7195));
assign g21760 = ((~g20198))|((~g6369));
assign g15804 = ((~g11660))|((~g12392));
assign g19296 = ((~II25624))|((~II25625));
assign g29134 = ((~II38145));
assign II25840 = ((~g17802))|((~II25838));
assign g11054 = ((~II17969));
assign g21421 = (g15274&g20411);
assign g22914 = ((~g21874))|((~g21871))|((~g21868));
assign g18617 = ((~g16094)&(~g14606));
assign g12249 = ((~g10510)&(~g10568)&(~g10613));
assign g13364 = ((~II20451));
assign g17442 = ((~II23530));
assign g25258 = ((~g24846)&(~g23741));
assign g10517 = (g3650&g5078);
assign g5904 = ((~g1224));
assign II15484 = ((~g3249));
assign g16291 = (g5855&g11931);
assign g12899 = ((~g8483)&(~g8498)&(~g8511));
assign g30690 = ((~g13489)&(~g30352));
assign II19289 = ((~g10653));
assign II20462 = ((~g10825));
assign g28630 = ((~g28118));
assign g13088 = ((~g9534))|((~g6912));
assign II37005 = ((~g28077));
assign g24708 = ((~g23854)&(~g22727));
assign g24299 = ((~II31571));
assign II36656 = ((~g27311));
assign g12025 = ((~g11355));
assign g22026 = ((~g21083)&(~g18407));
assign g25989 = ((~II33819));
assign II40571 = ((~g30588))|((~g30632));
assign g29324 = ((~g28718)&(~g19124));
assign g22380 = ((~g20833));
assign g4357 = ((~g729));
assign g24028 = ((~g22922))|((~g14135));
assign g29651 = ((~II39071));
assign g13510 = ((~g12565))|((~g3254));
assign II19826 = ((~g10252));
assign II37481 = ((~g27763));
assign g30918 = (g30780&g22296);
assign g23329 = ((~g22165)&(~g10133));
assign g20647 = (g5888&g19075);
assign g19258 = ((~II25525));
assign g22543 = ((~II29093));
assign II31820 = ((~g23844));
assign g13440 = ((~II20619));
assign g28194 = ((~II36860));
assign g23575 = ((~II30651));
assign II36618 = ((~g27300));
assign g30874 = ((~II40874));
assign II35551 = ((~g27075));
assign g25703 = ((~II33529));
assign g25569 = ((~g24708)&(~g24490));
assign g30911 = ((~II40985));
assign g12035 = ((~g10203)&(~g10289)&(~g10367));
assign g21359 = ((~II27900));
assign g26649 = ((~g25827));
assign g22668 = ((~g16075))|((~g21271));
assign II18551 = ((~g8824));
assign II21841 = ((~g13109));
assign g28124 = ((~II36797));
assign g26555 = ((~g25507));
assign g24081 = ((~g22852))|((~g14102));
assign g5833 = ((~g2133));
assign II14590 = ((~g1148));
assign II20682 = ((~g11659));
assign II32133 = ((~g24214));
assign g27992 = ((~II36473));
assign g19783 = ((~II26220));
assign g9745 = (g3722&g3981);
assign g28247 = ((~II36990));
assign g26086 = ((~II33984));
assign g23025 = ((~g21762)&(~g21124));
assign g19640 = ((~g16940));
assign g7819 = ((~g479));
assign II32198 = ((~g24250));
assign g27588 = ((~g26947)&(~g24742));
assign g23830 = (g22958&g9670);
assign g19689 = ((~II26112));
assign g16162 = (g5597&g13234);
assign g29650 = ((~II39068));
assign g29971 = (g29763&g13861);
assign g30906 = ((~II40970));
assign II26535 = ((~g18218));
assign g27951 = (g4438&g27459);
assign g13178 = ((~g9384));
assign g30566 = ((~g14327)&(~g30398));
assign g30247 = ((~g16112)&(~g30080));
assign g25992 = ((~II33828));
assign g27910 = ((~II36367));
assign II23983 = ((~g9216))|((~II23981));
assign g25442 = ((~II33265));
assign g4626 = ((~g735));
assign II37662 = ((~g28447));
assign II14637 = ((~g1849));
assign II20049 = ((~g10185))|((~II20048));
assign II16942 = ((~g7195));
assign g20242 = ((~g16852));
assign g24585 = (g2147&g23473);
assign g19322 = ((~g16636));
assign g25962 = ((~g24591)&(~g23496));
assign g23858 = ((~g23025)&(~g18554)&(~g4632));
assign II23733 = ((~g14831));
assign g8286 = ((~g3461));
assign g11398 = ((~II18356));
assign g5190 = ((~g2101));
assign g13479 = (g6017&g12196);
assign g22537 = ((~II29087));
assign II21688 = ((~g11699));
assign g12228 = ((~II19404));
assign g25056 = ((~g24242)&(~g17065));
assign g28637 = ((~g28192)&(~g17100));
assign g27273 = ((~g27001)&(~g26307));
assign II25210 = ((~g18986));
assign g25700 = ((~II33526));
assign g26746 = ((~II34845));
assign g8459 = (g6838&g2297);
assign g10486 = ((~g7957));
assign II30101 = ((~g22734));
assign g22069 = ((~g19477))|((~g21253))|((~g19522));
assign II40982 = ((~g30802));
assign g19319 = ((~g16633));
assign g4016 = ((~g417));
assign g25483 = (g24481&g20421);
assign g11123 = ((~II18037));
assign g30095 = (g29857&g11265);
assign g6518 = ((~II14775));
assign g24326 = ((~II31652));
assign g24258 = (g19481)|(g22404);
assign g18590 = ((~g16439)&(~g7522));
assign II27293 = ((~g19335));
assign II32478 = ((~g17927))|((~g24065));
assign g20505 = ((~g18371));
assign II29503 = ((~g21016));
assign g6020 = ((~g1573));
assign g26187 = ((~II34091));
assign g23864 = (g18297&g23057);
assign gbuf21 = (g3117);
assign g6047 = ((~g2285));
assign g28276 = ((~II37077));
assign g17774 = (g4696&g15429);
assign g20423 = ((~g17658));
assign II17881 = ((~g7976));
assign g29403 = ((~g28836)&(~g28383));
assign g26424 = (g5110&g25752);
assign g5411 = ((~II13947));
assign g29768 = ((~g29469)&(~g19146));
assign g30551 = ((~II40233));
assign g22093 = ((~g19500))|((~g21261))|((~g19532));
assign II24285 = ((~g15992));
assign g11011 = ((~II17922));
assign g17520 = ((~II23608));
assign g22984 = (g16840&g21400);
assign g28424 = (g17741&g28153);
assign g17015 = (g7996&g15390);
assign g24290 = ((~II31544));
assign II29981 = ((~g22702));
assign g24269 = ((~II31481));
assign II18590 = ((~g8793));
assign II18710 = ((~g8827));
assign g29814 = (g29728&g22266);
assign g4369 = ((~g852));
assign g16842 = ((~II22810));
assign g16643 = ((~g15904)&(~g14642)&(~g15859));
assign II21160 = ((~g12538));
assign g28915 = (g28619&g9323);
assign g20694 = ((~II27285));
assign g19521 = (g15080)|(g16781);
assign g22516 = (g20885&g17442);
assign g29989 = (g29893&g8391);
assign g29967 = (g29754&g12066);
assign g24317 = ((~II31625));
assign II28100 = ((~g19987));
assign g19984 = ((~g17197))|((~g780));
assign g7888 = ((~g1858));
assign g14177 = ((~g12920));
assign II13956 = ((~g1742));
assign II37781 = ((~g28595));
assign g18166 = ((~II24171));
assign II31637 = ((~g23663));
assign g11683 = ((~g9534))|((~g3366));
assign g30549 = ((~II40227));
assign II35723 = ((~g27168));
assign g13933 = (g7632&g12853);
assign g8973 = ((~II16283));
assign g10883 = ((~II17746));
assign g4523 = ((~g1397));
assign g16064 = ((~g12808));
assign II34863 = ((~g26576));
assign II20299 = ((~g10800));
assign g29678 = ((~g29545)&(~g29323));
assign II25222 = ((~g19011));
assign g16153 = (g5592&g13229);
assign g25472 = ((~II33300));
assign II38208 = ((~g28839));
assign g25698 = ((~g24600));
assign g10601 = ((~II17527));
assign g30067 = ((~g29818)&(~g29820));
assign g21301 = (g9453&g20289);
assign g11711 = ((~g9138)&(~g9143)&(~g9145));
assign II16793 = ((~g7265));
assign II37617 = ((~g28607));
assign g21975 = ((~g21245)&(~g21259));
assign g23179 = ((~II29990));
assign g7700 = ((~g3096));
assign g20735 = ((~II27324));
assign g11312 = ((~II18262));
assign II26401 = ((~g17012));
assign II22972 = ((~g9174))|((~g13962));
assign g11516 = ((~II18524));
assign g16394 = (g1675&g12054);
assign g30597 = ((~g6119)&(~g30412)&(~g25341));
assign g29486 = (g21544&g29291);
assign g28317 = ((~II37200));
assign g7865 = ((~g2554));
assign g12461 = ((~II19645));
assign g4902 = ((~g721));
assign II33837 = ((~g25723));
assign g19708 = (g1319&g18841);
assign g4668 = ((~g1418));
assign g19596 = ((~II26028));
assign g19865 = ((~g16607))|((~g9636));
assign g16178 = (g2372&g11846);
assign g20400 = ((~g17567));
assign g24162 = ((~g22552));
assign g30695 = ((~g13515)&(~g30374));
assign g8522 = (g6519&g957);
assign II36939 = ((~g28095));
assign g11497 = ((~II18467));
assign II23923 = ((~g13563));
assign g22134 = ((~g21803))|((~g21809));
assign g13863 = ((~II20959));
assign g6979 = ((~II14874));
assign II40679 = ((~g30641));
assign II23123 = ((~g9374))|((~g13866));
assign g19241 = (g16867&g14158&g14071);
assign II18184 = ((~g5837));
assign g9666 = ((~II16759));
assign g4281 = ((~g1792));
assign g9143 = (g7265&g7812);
assign g4360 = ((~g819));
assign g5685 = ((~g988));
assign g23232 = ((~II30149));
assign g22487 = ((~II29033));
assign g26335 = (g25907&g9666);
assign g9303 = ((~II16538));
assign g19109 = (g13724&g16360&II25300);
assign g4055 = ((~g1529));
assign g16299 = (g5860&g11941);
assign g19823 = (g4711&g17782);
assign g18245 = (g5283&g15744);
assign g15526 = (g5033&g13232);
assign g29432 = ((~II38677));
assign g4754 = ((~g713));
assign g15411 = (g4787&g13209);
assign g9229 = ((~II16499));
assign g13354 = ((~g8183)&(~g8045)&(~g11190)&(~g7880));
assign g15492 = ((~g12318));
assign g15382 = ((~II21644));
assign g8230 = ((~g1530));
assign g28768 = ((~II37729));
assign II25571 = ((~g740))|((~g18286));
assign g21802 = (g20147)|(g20119)|(II28323);
assign II36888 = ((~g27988));
assign g9880 = ((~II16876));
assign g25844 = ((~II33686));
assign g10641 = (g7303&g2679);
assign g28133 = ((~g27550));
assign II13538 = ((~g2870));
assign II29999 = ((~g22756));
assign g12119 = ((~g11475));
assign g28011 = ((~II36510));
assign g28332 = (g27883&g22331);
assign g20463 = ((~g17856));
assign g13289 = (g5647&g11141);
assign g10909 = ((~II17786));
assign g26151 = ((~g6068)&(~g24183)&(~g25335));
assign g12042 = ((~g11373));
assign g21401 = (g9507&g20397);
assign g19556 = ((~II25985));
assign g12597 = ((~g8752));
assign II40565 = ((~g30700));
assign g6042 = ((~II14519));
assign II38128 = ((~g28419));
assign g29889 = ((~g29684));
assign II24171 = ((~g16439));
assign g29519 = ((~II38885));
assign g19928 = (g2740&g18964);
assign II25264 = ((~g17151));
assign g23258 = ((~II30227));
assign g7858 = ((~g1164));
assign g12881 = ((~g8918));
assign g23169 = ((~II29960));
assign g21255 = ((~g20022)&(~g5963));
assign II35814 = ((~g27125));
assign II30844 = ((~g22102));
assign II40251 = ((~g30463));
assign g13519 = ((~g13228));
assign II33232 = ((~g24863));
assign g27376 = ((~II35698));
assign g25392 = (g24700&g18400);
assign g12295 = ((~g8478));
assign g27501 = ((~g26763)&(~g24436));
assign g13029 = ((~g9676))|((~g7162));
assign II30056 = ((~g22589));
assign g26040 = (g25745&g19533);
assign gbuf32 = (g282);
assign gbuf48 = (g397);
assign g16476 = ((~II22530));
assign II32112 = ((~g24207));
assign II16664 = ((~g7265));
assign g10623 = (g3650&g5249);
assign g9730 = ((~II16779));
assign II23424 = ((~g15826));
assign g7739 = ((~g1700));
assign g16480 = ((~II22542));
assign g18483 = ((~g14573));
assign II37880 = ((~g28529));
assign II29418 = ((~g20982));
assign g5692 = ((~g1501));
assign II22575 = ((~g15092));
assign II29197 = ((~g20903));
assign g18088 = (g5150&g15667);
assign gbuf28 = (g450);
assign II30547 = ((~g23093));
assign II16279 = ((~g5419));
assign II31703 = ((~g23861));
assign II38080 = ((~g28358));
assign g11704 = ((~g9822))|((~g3678));
assign g11243 = ((~II18169));
assign II16131 = ((~g5408));
assign g18857 = ((~g15343));
assign g10412 = (g3834&g4870);
assign g21757 = (g3866&g20554);
assign II34086 = ((~g25215));
assign II22618 = ((~g14630));
assign gbuf87 = (g1037);
assign g5755 = ((~g240));
assign II22611 = ((~g15055));
assign g21893 = ((~g13541)&(~g19328));
assign g15887 = ((~g12611))|((~g6369));
assign g14711 = ((~II21274));
assign g22150 = ((~g21420)&(~g19746));
assign g16046 = (g5618&g11761);
assign g20296 = ((~g17272));
assign g28998 = ((~II37961));
assign g28699 = ((~II37644));
assign g5266 = ((~g2523));
assign g30763 = (g30597&g22386);
assign II39398 = ((~g29664));
assign g21004 = ((~g19826)&(~g17874));
assign II39674 = ((~g30072));
assign g11846 = ((~g11056));
assign II20541 = ((~g11599));
assign g14991 = ((~g12262));
assign g23058 = ((~g16999)&(~g21112));
assign g16053 = (g297&g11770);
assign g12471 = ((~II19657));
assign II14990 = ((~g2697));
assign II27029 = ((~g19176));
assign II14587 = ((~g1085));
assign II15602 = ((~g6783));
assign II23527 = ((~g15858));
assign g10573 = (g5512&g5173);
assign g11252 = ((~II18178));
assign II24362 = ((~g6157))|((~II24361));
assign g18307 = ((~g14298));
assign g24504 = ((~g23770)&(~g23818));
assign II34096 = ((~g25218));
assign II17235 = ((~g3900));
assign g26878 = ((~g26482)&(~g5680));
assign g15435 = (g4702&g12801);
assign g27695 = ((~II36096));
assign II27749 = ((~g19954));
assign II34220 = ((~g25248));
assign g22227 = ((~g21658)&(~g19953));
assign II35791 = ((~g26779));
assign gbuf154 = (g1950);
assign g23438 = ((~II30467));
assign g4942 = ((~g1422));
assign II29939 = ((~g22518));
assign II36371 = ((~g27674));
assign g30671 = ((~g16391)&(~g30486));
assign g3461 = ((~g992));
assign g13452 = ((~II20655));
assign g29467 = (g29340&g19467);
assign g20892 = ((~g19627)&(~g17448));
assign g20310 = ((~g16850)&(~g13654));
assign II13143 = ((~g39));
assign g27771 = ((~g27578)&(~g27115));
assign II39026 = ((~g29510));
assign g25729 = ((~II33558));
assign g30770 = ((~II40568));
assign II22414 = ((~g1206));
assign g17419 = ((~II23507));
assign II15350 = ((~g2549));
assign g12657 = ((~II19777));
assign II25365 = ((~g18707));
assign g24036 = ((~g22852))|((~g14467));
assign g27364 = (g1435&g26855);
assign g25173 = ((~II32997));
assign II37871 = ((~g28556));
assign g25523 = ((~g20842)&(~g24429));
assign g20452 = ((~g17782));
assign g16676 = ((~II22718));
assign g28685 = ((~II37602));
assign g9787 = ((~II16835));
assign g25761 = ((~g25112)&(~g6305));
assign gbuf140 = (g1748);
assign g22761 = ((~II29503));
assign g13121 = ((~g9968))|((~g7426));
assign g13317 = ((~II20376));
assign g29298 = ((~II38437));
assign g23248 = ((~II30197));
assign g14347 = ((~g12079));
assign g13035 = ((~g9534))|((~g6912));
assign g21781 = ((~g20255))|((~g7085));
assign gbuf59 = (g566);
assign g5394 = ((~g3054));
assign g28512 = (g26481)|(g27738);
assign g19727 = (g4329&g17557);
assign g15074 = ((~g11962));
assign g4955 = ((~g1905));
assign II29468 = ((~g21003));
assign II14865 = ((~g1237));
assign g26193 = ((~II34105));
assign g24057 = ((~g22922))|((~g14626));
assign g15678 = ((~g12382));
assign g4301 = ((~g2233));
assign g26505 = ((~II34473));
assign g12821 = ((~g8863));
assign g28232 = ((~II36945));
assign II34277 = ((~g25257));
assign II24647 = ((~g14385))|((~II24646));
assign II36072 = ((~g27480));
assign g21874 = ((~g18561))|((~g19233))|((~g19244));
assign g26347 = (g25915&g9730);
assign g10915 = ((~II17798));
assign II21252 = ((~g11644));
assign II37752 = ((~g28512));
assign g14546 = ((~g12213));
assign g10388 = (g3618&g4818);
assign g21670 = (g3554&g20505);
assign g24487 = ((~g23666)&(~g23709));
assign II17756 = ((~g7192));
assign g15588 = ((~II21844));
assign g5728 = (g1024&g1040);
assign g5320 = ((~g2793));
assign g28079 = (g27599&g10127);
assign g19945 = ((~II26401));
assign II29579 = ((~g21043));
assign g16418 = (g5959&g12084);
assign g11567 = ((~II18677));
assign g18930 = ((~g15612));
assign g26852 = ((~II35007));
assign II33347 = ((~g24438));
assign II28178 = ((~g20067));
assign II19997 = (g9391&g9326&g9264&g9216);
assign II26612 = ((~g17645));
assign II18990 = ((~g9183));
assign g24856 = ((~II32506));
assign II37146 = ((~g28108));
assign II39237 = ((~g29690));
assign g23678 = ((~II30832));
assign g4836 = ((~g2092));
assign II40495 = ((~g30680));
assign g8770 = ((~II15964));
assign g30678 = ((~g16427)&(~g30502));
assign II35394 = ((~g26183));
assign g19012 = ((~II25099));
assign g26182 = ((~II34086));
assign II23591 = ((~g14885));
assign g28152 = ((~g27391));
assign g16599 = ((~g14546));
assign g24757 = (g1358&g24110);
assign II30377 = ((~g22802));
assign g24773 = (g9711&g24125);
assign g19768 = (g17815&g16054);
assign II33790 = ((~g25103));
assign g7910 = ((~g474));
assign II22999 = ((~g9187))|((~II22998));
assign g13907 = ((~g12781));
assign g16140 = (g5705&g11825);
assign g12543 = ((~II19711));
assign g20430 = ((~g17682));
assign g16414 = (g5955&g12076);
assign g20411 = ((~g17607));
assign II20417 = ((~g10933));
assign g24574 = (g23441&g18240&g23100);
assign g23896 = ((~II31162));
assign g19194 = (g18492)|(g17830);
assign g19577 = ((~g16881));
assign g15609 = ((~II21865));
assign g20040 = ((~II26476));
assign g27464 = ((~g27178)&(~g25975));
assign g15201 = ((~II21491));
assign g8726 = ((~II15932));
assign g8093 = ((~g2972));
assign g25714 = ((~II33542));
assign g18222 = (g5257&g15731);
assign g5717 = ((~g793));
assign g29474 = (g21508&g29271);
assign II26661 = (g18679&g18699&g16201);
assign g11888 = ((~g11021));
assign g24449 = ((~g23694))|((~g3462));
assign g29570 = ((~g28709)&(~g29175));
assign II32347 = ((~g24002))|((~II32345));
assign g4139 = ((~g867));
assign II18323 = ((~g6369));
assign II40450 = ((~g30592));
assign g12363 = ((~II19523));
assign g11341 = ((~II18295));
assign g7580 = ((~g2568));
assign g17218 = ((~g15933)&(~g14669));
assign g30297 = ((~g13490)&(~g29994));
assign II36667 = ((~g27551))|((~II36666));
assign g23038 = ((~g21566));
assign g19482 = ((~g17194));
assign II23008 = ((~g9203))|((~g13926));
assign g23414 = (g21569&g22421);
assign g24491 = ((~g15247)&(~g23735));
assign g23823 = ((~g23009)&(~g18490)&(~g4456));
assign g17576 = (g4348&g15248);
assign g12513 = ((~g8651));
assign g22597 = (g21921&g12708);
assign g18815 = ((~g15161));
assign II31583 = ((~g23783));
assign g25246 = ((~g24810)&(~g23637));
assign gbuf169 = (g2214);
assign g5957 = ((~g273));
assign g9423 = ((~g5428));
assign II27092 = ((~g19174));
assign g11417 = ((~II18381));
assign II17789 = ((~g7388));
assign g7333 = ((~g2358));
assign II29354 = ((~g20964));
assign g26671 = ((~g25226)&(~g10238));
assign g11294 = ((~II18244));
assign g10767 = ((~g6294));
assign g8792 = ((~II15992));
assign g30988 = ((~II41138));
assign g6161 = ((~g1210));
assign g7837 = ((~g3044));
assign II40614 = ((~g30709));
assign II33501 = ((~g25057));
assign g30101 = (g29857&g11341);
assign g10796 = ((~II17641));
assign g11920 = ((~g11182));
assign g22629 = ((~II29229));
assign g24964 = (g7595&g24251);
assign g23477 = ((~g22906)&(~g21758));
assign g25212 = ((~g24751)&(~g23559));
assign g4976 = ((~g2113));
assign g13133 = ((~g9968))|((~g7488));
assign gbuf202 = (g2638);
assign g7642 = ((~g3125));
assign g20966 = ((~g19765)&(~g17734));
assign g25278 = (g24668&g8719);
assign g27391 = ((~II35731));
assign g10848 = ((~g5801));
assign g23273 = ((~II30272));
assign g22995 = ((~g21441));
assign II16206 = ((~g6448));
assign g29760 = ((~g16411)&(~g29624));
assign g15425 = (g4832&g13212);
assign II19901 = ((~g10746));
assign g25404 = ((~g24771));
assign II38613 = ((~g28886));
assign g25631 = ((~g24717)&(~g24497));
assign g19653 = (g4095&g17430);
assign g25457 = (g6163&g24784);
assign g19456 = ((~II25898))|((~II25899));
assign II24624 = ((~g6136))|((~g14252));
assign g23237 = ((~II30164));
assign II29506 = ((~g21017));
assign g12755 = ((~g11431)&(~g8339)&(~g8394));
assign g13352 = ((~g10419));
assign g18212 = ((~II24214))|((~II24215));
assign g28971 = (g28630&g9501);
assign g26771 = (g24912&g26508&g13614);
assign g22130 = ((~g21393)&(~g19711));
assign g17926 = (g4936&g15553);
assign g29187 = ((~g28854)&(~g28416));
assign g21028 = ((~g19863)&(~g15591));
assign g5113 = ((~g2519));
assign g8028 = ((~g3078));
assign g27897 = ((~g6087)&(~g27632)&(~g25349));
assign g15596 = ((~II21852));
assign g15544 = ((~g12340));
assign g13260 = ((~g10067));
assign g26249 = ((~II34201));
assign g26705 = ((~II34722));
assign g19657 = ((~II26085));
assign II31053 = ((~g22163));
assign g29576 = ((~g28713)&(~g29183));
assign II16741 = ((~g6062));
assign g21990 = (g291&g21187);
assign II41117 = ((~g30977));
assign g24748 = (g672&g24101);
assign II14056 = ((~g1880));
assign g16859 = (g15762&g8662);
assign g28227 = ((~II36930));
assign g22263 = ((~g21723)&(~g20021));
assign g30289 = ((~g16458)&(~g29985));
assign g29285 = ((~g28804));
assign g22172 = ((~g21455)&(~g19790));
assign g8153 = ((~g1527));
assign g20045 = ((~II26481));
assign g23132 = ((~g17155)&(~g21209));
assign g22049 = ((~g21315)&(~g19576));
assign II33268 = ((~g24925));
assign II40161 = ((~g30439));
assign g29158 = ((~II38217));
assign II33819 = ((~g25707));
assign II36972 = ((~g28052));
assign g21210 = (g20242&g12415);
assign II16325 = ((~g6052));
assign g30754 = (g30614&g22313);
assign g26550 = ((~g25493));
assign II27766 = ((~g19984));
assign II29313 = ((~g20948));
assign g29167 = ((~g28841)&(~g28396));
assign g30591 = ((~II40317));
assign g20001 = (g5355&g18450);
assign g20349 = ((~g17405));
assign g27599 = ((~g27147));
assign g27238 = ((~II35551));
assign II29058 = ((~g20703));
assign g30669 = ((~g16383)&(~g30481));
assign g15284 = ((~II21560));
assign g25422 = ((~g24958));
assign g23239 = ((~II30170));
assign g8538 = (g6783&g1570);
assign g26351 = (g4865&g25623);
assign II16857 = ((~g7053));
assign g25076 = ((~g23409)&(~g22187));
assign II16482 = ((~g6000));
assign g19200 = (g18346)|(g18424);
assign g29343 = ((~g28338)&(~g28724));
assign g12219 = ((~g8414));
assign g20884 = ((~g5394)&(~g19830));
assign g16430 = (g5974&g12116);
assign g29708 = ((~II39168));
assign g22097 = ((~g21355)&(~g19649));
assign g13426 = ((~II20577));
assign II26846 = ((~g17229));
assign g17490 = ((~II23578));
assign g23435 = ((~g23120));
assign II36081 = ((~g27497));
assign g7478 = ((~g1138));
assign II31302 = ((~g22284));
assign g29039 = ((~g28322)&(~g13500));
assign g25944 = ((~g24542)&(~g24552));
assign II14191 = ((~g2400));
assign II27658 = ((~g20526));
assign g23151 = ((~II29906));
assign g24660 = ((~g2574))|((~g23402));
assign g27110 = (g5298&g26485);
assign g18678 = ((~g13625)&(~g11771));
assign II20379 = ((~g11213));
assign g10567 = (g6945&g5159);
assign g29307 = ((~II38456));
assign II39926 = ((~g30296));
assign II25219 = ((~g19009));
assign g29275 = ((~g28779));
assign g10116 = (g6519&g4360);
assign g23319 = (g14493)|(g22385);
assign II30224 = ((~g22795));
assign g23470 = ((~g22188));
assign g22242 = ((~g21687)&(~g19983));
assign g21336 = (g9203&g20332);
assign II16850 = ((~g3618));
assign II23287 = ((~g13741));
assign g30712 = ((~II40426));
assign g30970 = ((~g30917)&(~g30921)&(~g30953));
assign g23014 = ((~g16939)&(~g21077));
assign g28063 = ((~II36636));
assign g13244 = ((~g10004));
assign g24555 = ((~g23912)&(~g22798));
assign g17754 = (g4662&g15418);
assign g16103 = (g5621&g11796);
assign g22826 = ((~g16113)&(~g20904));
assign g15308 = ((~II21577));
assign II39828 = ((~g30269));
assign g21391 = (g15188&g20386);
assign II15562 = ((~g5778));
assign g10093 = (g7426&g4315);
assign g5911 = ((~g1889));
assign II24566 = ((~g14472))|((~II24565));
assign g27158 = ((~II35355));
assign g19281 = (g17171)|(g17150)|(II25588);
assign g12959 = ((~g8513)&(~g8528)&(~g8543));
assign g26575 = ((~g13845)&(~g25295));
assign II25402 = ((~g18821));
assign g23938 = ((~g22852))|((~g14028));
assign g24885 = (g18374&g23839);
assign g4089 = ((~g2836));
assign II29569 = ((~g21040));
assign g13224 = ((~g9819));
assign II29043 = ((~g21748));
assign II39690 = ((~g30035))|((~II39689));
assign g10590 = (g7265&g5204);
assign II26558 = (g14776&g18670&g18720);
assign g13833 = (g7919&g12009);
assign g11303 = ((~II18253));
assign II35020 = ((~g26110))|((~g26099));
assign g17746 = ((~II23821));
assign II29924 = ((~g23094));
assign g5404 = ((~II13928));
assign g22872 = ((~II29672));
assign II31517 = ((~g23641));
assign II40447 = ((~g30587));
assign g22062 = (g21135&g21118&g21106&II28609);
assign g13099 = ((~g9534))|((~g6912));
assign II39080 = ((~g29568));
assign g20361 = ((~g17430));
assign g12425 = ((~II19573));
assign g25051 = ((~g23803))|((~g7265));
assign g15566 = ((~II21822));
assign II37035 = ((~g28017));
assign g15423 = (g4827&g13210);
assign g8285 = ((~g3365));
assign g24152 = ((~g22533));
assign II33448 = ((~g25050));
assign g11003 = ((~II17910));
assign g25410 = ((~g24723));
assign g21742 = ((~g19919));
assign g30533 = ((~II40179));
assign II25374 = ((~g18726));
assign g12791 = ((~II19852));
assign g15357 = ((~II21626));
assign g22418 = ((~II28962));
assign g19022 = ((~II25129));
assign g18918 = ((~II24950));
assign g29338 = (g29060&g29042);
assign II37014 = ((~g28097));
assign g30339 = ((~II39848));
assign II40670 = ((~g30638));
assign g25420 = ((~II33246));
assign II19736 = ((~g9184));
assign g5844 = ((~g2377));
assign g26060 = (g25943&g21108);
assign gbuf80 = (g967);
assign g25882 = ((~g4632)&(~g25082)&(~g18502)&(~g16113));
assign g28993 = ((~II37956));
assign g22113 = ((~g21371)&(~g19671));
assign II38812 = ((~g15904))|((~II38810));
assign g17395 = (g6177&g15034);
assign g3254 = ((~II13158));
assign g7015 = ((~II14885));
assign g21765 = ((~g20228))|((~g6783));
assign g27066 = ((~g26024)&(~g20665));
assign II19711 = ((~g10230));
assign II23057 = ((~g13982))|((~II23055));
assign g18651 = (g14863&g15065&g16266&g13819);
assign II17804 = ((~g8031));
assign g19743 = (g1346&g18858);
assign g8351 = ((~II15553));
assign II40059 = ((~g30259));
assign g17919 = ((~II23967))|((~II23968));
assign g29068 = ((~g9326))|((~g28567));
assign II33822 = ((~g25770));
assign g28672 = (g27950&g13859);
assign II21586 = ((~g13054));
assign g26008 = ((~II33876));
assign g21147 = ((~g20135)&(~g20158)&(~g20188));
assign g24071 = ((~g22852))|((~g14201));
assign g22991 = ((~g21429));
assign g26382 = (g25915&g9812);
assign II18554 = ((~g8866));
assign g21912 = (g19327&g13011);
assign II39391 = ((~g29769))|((~g15971));
assign g12001 = ((~g11315));
assign g24534 = ((~g15561)&(~g23893));
assign II36337 = ((~g27628));
assign g10198 = (g6643&g571);
assign g4693 = ((~g2084));
assign g11082 = ((~II17992));
assign g28031 = ((~II36554));
assign g30600 = ((~II40326));
assign g17697 = (g4555&g15363);
assign g15225 = ((~II21508));
assign II17527 = ((~g3900));
assign g23785 = ((~II30997));
assign g18205 = ((~g14467));
assign g23418 = ((~g17794)&(~g22690));
assign g11553 = ((~II18635));
assign g18463 = ((~g14408));
assign g13239 = ((~g9933));
assign g27313 = ((~g27055)&(~g26400));
assign g29621 = ((~g14059)&(~g29263));
assign II15299 = ((~g1168));
assign g27472 = ((~II35814));
assign II33636 = ((~g24525));
assign II32266 = ((~g17903))|((~II32265));
assign g19223 = (g18195)|(g18290);
assign g27176 = ((~II35383));
assign II24718 = ((~g9941))|((~II24716));
assign g27810 = ((~g27632)&(~g1215));
assign II27221 = ((~g19180));
assign g25943 = ((~g24541)&(~g24550));
assign II23199 = ((~g9569))|((~II23198));
assign g5167 = ((~g1410));
assign g19094 = (g18679&g14849&g16254&g13756);
assign g30664 = ((~g16358)&(~g30473));
assign g13419 = ((~II20556));
assign II14238 = ((~g2406));
assign g16487 = ((~II22563));
assign II29392 = ((~g20975));
assign II29151 = ((~g20893));
assign g17130 = ((~g13541));
assign g18913 = ((~II24943));
assign g24000 = ((~II31232));
assign g25273 = ((~g24907)&(~g23904));
assign g24516 = ((~g23820)&(~g22700));
assign II33627 = ((~g25059));
assign II32401 = ((~g17927))|((~II32400));
assign g3251 = ((~II13149));
assign g29645 = ((~II39053));
assign g21228 = ((~g19388)&(~g17118));
assign g27179 = ((~g26082)&(~g25356));
assign g23566 = ((~II30632));
assign II34824 = ((~g26282));
assign g13414 = ((~II20541));
assign g28427 = (g26092&g28154);
assign g10445 = (g6945&g1285);
assign II38056 = ((~g28351));
assign g5898 = ((~g762));
assign II25528 = ((~g18942));
assign g30237 = ((~g30032));
assign g10285 = (g6486&g4606);
assign II28767 = ((~g13552))|((~II28765));
assign g16110 = (g516&g11804);
assign II29262 = ((~g20926));
assign g23820 = (g3013&g23036);
assign g17893 = ((~g14165));
assign g6304 = ((~g1672));
assign g10859 = ((~II17712));
assign g17028 = (g7604&g15458);
assign II31014 = ((~g22152));
assign g20107 = (g18415&g3173);
assign g12945 = (II19996&II19997);
assign II21277 = ((~g12430));
assign g30654 = ((~g16299)&(~g30457));
assign g24046 = ((~g22922))|((~g14637));
assign g12951 = ((~g8993));
assign g29978 = ((~II39472));
assign II31270 = ((~g22247));
assign II27422 = ((~g19431));
assign g20584 = ((~II27077));
assign g22674 = (g14092&g21537);
assign II24213 = ((~g14033))|((~g9711));
assign II30826 = ((~g22097));
assign II30651 = ((~g22041));
assign g17842 = ((~g13936));
assign g24250 = ((~g17135)&(~g22358));
assign g25271 = ((~g24901)&(~g18047));
assign g23973 = ((~g22812))|((~g14450));
assign g23747 = (g18025&g23016);
assign g20112 = (g16749&g3132);
assign g27755 = ((~g27448)&(~g26986));
assign g18772 = ((~g15003));
assign II39086 = ((~g29497));
assign g16171 = ((~g10952)&(~g6188)&(~g12524));
assign g26399 = ((~g16571))|((~g25186));
assign II35744 = ((~g26906));
assign g21438 = (g9649&g20422);
assign II16939 = ((~g3650));
assign g29697 = ((~II39145));
assign g21039 = ((~g19879)&(~g18035));
assign II18169 = ((~g7195));
assign g25724 = ((~II33554));
assign II36769 = ((~g27340));
assign g29920 = ((~g24723)&(~g29739));
assign g5015 = ((~g2788));
assign g21866 = ((~g18363))|((~g19212))|((~g19222));
assign g12521 = ((~g8659));
assign g21606 = ((~II28137));
assign g10931 = ((~II17816));
assign II23942 = ((~g13946))|((~II23941));
assign gbuf132 = (g1667);
assign g13496 = (g6032&g12246);
assign g5640 = ((~g3170));
assign g20500 = ((~g18278));
assign g14618 = ((~g11844));
assign II33577 = ((~g24462));
assign II32934 = ((~g25123));
assign g13143 = ((~g8636)&(~g8654)&(~g8666));
assign II22925 = ((~g15118))|((~II22924));
assign g29476 = (g21544&g29274);
assign g15322 = ((~g12239));
assign gbuf149 = (g1925);
assign II25096 = ((~g15161));
assign g23719 = ((~II30891));
assign g11747 = ((~g10898));
assign g23260 = ((~II30233));
assign II36975 = ((~g28032));
assign II39906 = ((~g30290));
assign II40134 = ((~g30480));
assign II35022 = ((~g26099))|((~II35020));
assign II30308 = ((~g22725));
assign g25780 = ((~II33617));
assign g20545 = ((~g18519));
assign g15623 = (g5185&g13260);
assign g24228 = ((~g17028)&(~g22285));
assign g9161 = ((~g5852));
assign II39463 = ((~g29933));
assign g30769 = ((~II40565));
assign g27734 = (g27538&g16814);
assign g4862 = ((~g2418));
assign g28368 = ((~g15770)&(~g28123));
assign g12129 = (g7872&g8788);
assign II38692 = ((~g29317));
assign g22222 = ((~g21935));
assign g8650 = (g7053&g7224);
assign g25120 = ((~g23901));
assign II31159 = ((~g22192));
assign g27187 = (g16594&g26516&g13626);
assign II15574 = ((~g6838));
assign g18890 = ((~II24916));
assign II21259 = ((~g11630));
assign g28445 = (g26121&g28164);
assign gbuf58 = (g574);
assign g15878 = ((~g13375))|((~g12392));
assign g13100 = ((~g9534))|((~g6678));
assign II30480 = ((~g23014));
assign g28823 = ((~II37784));
assign II13677 = ((~g809));
assign II25839 = ((~g88))|((~II25838));
assign g8811 = ((~II16021));
assign g26653 = ((~g25844));
assign II22632 = ((~g15978))|((~II22630));
assign g21252 = (g19578&g14895);
assign II19615 = ((~g10789));
assign g30557 = ((~II40251));
assign II32210 = ((~g23539));
assign g23734 = (g17974&g23008);
assign g4869 = ((~g2513));
assign g25552 = (g7009&g25104);
assign g18079 = ((~II24092))|((~II24093));
assign g10966 = ((~II17857));
assign g30381 = ((~II39948));
assign II40922 = ((~g30748));
assign g23554 = (g8147&g22418);
assign g10211 = (g6713&g1119);
assign g4165 = ((~g1553));
assign g21061 = ((~g19911)&(~g18153));
assign II15238 = ((~g2963))|((~II15237));
assign g9733 = ((~II16782));
assign g13943 = (g2622&g12867);
assign g18780 = ((~g13674)&(~g11847));
assign g19690 = ((~II26115));
assign g20825 = ((~g19219))|((~g15959));
assign g11912 = ((~g9931)&(~g10064)&(~g10155));
assign g23906 = ((~g22812))|((~g13958));
assign g15176 = ((~g12142));
assign g3305 = ((~g305));
assign g4860 = ((~II13652));
assign g19632 = (g4035&g17405);
assign g11985 = ((~g11291));
assign g27486 = ((~II35834));
assign II26491 = (g18497)|(g18441)|(g18363);
assign II36636 = ((~g27305));
assign g13188 = ((~g9465));
assign g10409 = ((~II17363));
assign g10404 = (g7265&g4862);
assign g6030 = ((~II14499));
assign g28618 = ((~g27861));
assign g24836 = ((~g16309)&(~g24241));
assign g15704 = ((~II21952));
assign g19906 = (g14614&g14048&II26354);
assign g10398 = (g7230&g4839);
assign g7852 = ((~g2981));
assign g4260 = ((~g1391));
assign g5000 = ((~g2459));
assign II39803 = ((~g30308));
assign II20667 = ((~g13396));
assign g24369 = ((~II31781));
assign g18841 = ((~g15265));
assign g3866 = ((~II13239));
assign II34967 = ((~g26553));
assign g15261 = ((~g12201));
assign g13094 = ((~g9822))|((~g7358));
assign II28896 = ((~g21246));
assign g13335 = (g5708&g11278);
assign g25350 = ((~II33182));
assign g8268 = ((~II15472));
assign g8933 = ((~II16225));
assign g30719 = ((~II40447));
assign II40182 = ((~g30332));
assign g8705 = (g3494&g7842);
assign II16450 = ((~g3834));
assign II34074 = ((~g25213));
assign g16491 = ((~II22575));
assign g20630 = ((~II27215));
assign II24667 = ((~g14559))|((~g9737));
assign g21619 = ((~II28148));
assign g20222 = (g18656&g18720&g13657&g16293);
assign g17168 = ((~g14041))|((~g13990));
assign g25222 = ((~g24768)&(~g23578));
assign g26669 = ((~g25360)&(~g17161));
assign II31035 = ((~g22941))|((~g14431));
assign g5301 = ((~g1964));
assign II16341 = ((~g7265));
assign g22287 = ((~g20735));
assign II33673 = ((~g24534));
assign II38091 = ((~g28362));
assign II37497 = ((~g27767));
assign g19135 = ((~g16739))|((~g16770));
assign II20506 = ((~g11189))|((~II20504));
assign II31553 = ((~g23501));
assign g23672 = (g4278&g22563);
assign g5596 = ((~II14052));
assign II23775 = ((~g15055));
assign g25499 = ((~II33327));
assign g16390 = (g982&g12041);
assign g14502 = ((~g12995));
assign g11903 = ((~g9912)&(~g10048)&(~g10122));
assign g3493 = ((~g996));
assign g27738 = ((~g25367))|((~g27415));
assign g17554 = (g4315&g15237);
assign II30140 = ((~g22623));
assign II34848 = ((~g26506));
assign II20607 = ((~g11990));
assign II18037 = ((~g7265));
assign g9954 = (g6838&g4188);
assign g5933 = ((~g873));
assign II30110 = ((~g22761));
assign II28330 = (g19099)|(g19094)|(g19089);
assign g26051 = (g70&g25296);
assign II27405 = ((~g19401));
assign g26268 = (g4509&g25507);
assign II34704 = ((~g26182));
assign II31037 = ((~g14431))|((~II31035));
assign g13655 = (g7540&g12518);
assign g27291 = ((~g27025)&(~g26350));
assign g9632 = (g6232&g3928);
assign II39641 = ((~g30057));
assign g4224 = ((~g429));
assign g17461 = (g6209&g15130);
assign g12009 = ((~II19195));
assign g13384 = ((~II20479));
assign II38085 = ((~g28360));
assign g4143 = ((~g1104));
assign II35479 = ((~g27171));
assign g22190 = (g16113)|(g20850);
assign g17354 = ((~II23442));
assign g23517 = ((~II30563));
assign g17499 = ((~g16292));
assign g24065 = ((~g22852))|((~g14286));
assign g26279 = (g25911&g9484);
assign g16824 = ((~g15658)&(~g12938));
assign g27699 = ((~II36108));
assign g12749 = ((~II19813));
assign II27101 = ((~g19220));
assign g13904 = (g7337&g12843);
assign g22156 = ((~II28693));
assign g29092 = ((~II38071));
assign g25506 = (g14263&g25095);
assign g26759 = (g26356&g19251);
assign II31091 = ((~g22173));
assign g23298 = ((~II30347));
assign II25830 = ((~g2138))|((~II25829));
assign g21772 = ((~g20255))|((~g7085));
assign g9910 = (g6713&g1098);
assign g8506 = (g6519&g948);
assign g22331 = ((~g20793));
assign g10130 = ((~II17106));
assign II15463 = ((~g3242));
assign g24345 = ((~II31709));
assign II35007 = ((~g26596));
assign II15317 = ((~g2842));
assign g29682 = ((~g29557)&(~g29336));
assign g21612 = ((~II28143));
assign g4674 = ((~g1511));
assign g17137 = ((~II23153))|((~II23154));
assign g21481 = (g9711&g20445);
assign g24375 = ((~II31799));
assign g12944 = ((~g8987));
assign g4124 = ((~g725));
assign g21739 = ((~g20507)&(~g18430));
assign II23412 = ((~g13482));
assign g26715 = ((~II34752));
assign II38238 = ((~g29119));
assign g6104 = ((~g1880));
assign g19348 = ((~II25741))|((~II25742));
assign g22584 = ((~II29148));
assign II40531 = ((~g30692));
assign g26830 = ((~II34961));
assign g27426 = ((~g27038))|((~g5512));
assign g10788 = ((~g7424));
assign g6053 = ((~II14538));
assign II30952 = ((~g22916))|((~g14309));
assign g17479 = ((~II23567));
assign II15184 = ((~g2975))|((~II15183));
assign g28847 = (g27850&g28609);
assign g6043 = ((~g1591));
assign g22280 = ((~g21749)&(~g20063));
assign II28800 = ((~g21316));
assign g25230 = ((~g24779)&(~g23598));
assign II18503 = ((~g8658));
assign g21790 = ((~g20228))|((~g6574));
assign II25771 = ((~g762))|((~g18436));
assign g24924 = (g24084&g18956);
assign g24907 = (g7466&g24220);
assign g10322 = (g7230&g4702);
assign II21491 = ((~g13038));
assign g11560 = ((~II18656));
assign g27081 = (g22108&g26638);
assign g16034 = ((~g12749));
assign g28293 = ((~II37128));
assign II39047 = ((~g29513));
assign g19050 = ((~II25213));
assign g24401 = ((~II31877));
assign II33431 = ((~g24450));
assign g24900 = ((~II32634))|((~II32635));
assign II36468 = ((~g27261));
assign II23364 = ((~g15805));
assign g29304 = ((~II38447));
assign g23802 = (g18142&g23032);
assign II17857 = ((~g6448));
assign II38345 = ((~g29109));
assign g19089 = (g14849&g18728&g16201&g16254);
assign II35044 = ((~g26145))|((~II35042));
assign g11861 = ((~g9766)&(~g9894)&(~g10013));
assign g30222 = (g30040&g9010);
assign g26494 = (g5315&g25865);
assign g10933 = ((~II17822));
assign II20743 = ((~g11621))|((~g13399));
assign II21942 = ((~g11724));
assign g29391 = ((~g29035));
assign g27722 = ((~g27252)&(~g10238));
assign II18113 = ((~g3997))|((~g8181));
assign g7542 = ((~g2883));
assign g9952 = (g3722&g4182);
assign g12552 = ((~II19722));
assign g28210 = ((~II36879));
assign g24319 = ((~II31631));
assign g17875 = (g4873&g15513);
assign II35099 = ((~g26672));
assign g17047 = (g7605&g15492);
assign II28057 = ((~g20067));
assign II14834 = ((~g1517));
assign g11641 = ((~II18827));
assign g11814 = (g1934&g8651);
assign g21690 = ((~g19098));
assign g5938 = ((~g1501));
assign II40946 = ((~g30726));
assign g23982 = ((~g22852))|((~g14580));
assign g14123 = ((~g11956));
assign II34752 = ((~g26220));
assign g30068 = ((~g29819)&(~g29821));
assign g21794 = ((~g19070)&(~g18617));
assign g23139 = (g5977&g21093);
assign g13571 = ((~II20791));
assign g5088 = ((~g1979));
assign II32976 = ((~g24588));
assign g5828 = (g1706&g1775);
assign II29323 = ((~g20951));
assign g4438 = ((~g2502));
assign II23788 = ((~g15901));
assign II37101 = ((~g27805));
assign g8408 = ((~II15610));
assign g16036 = ((~g6289)&(~g12467)&(~g10952));
assign g27180 = ((~II35389));
assign g20924 = ((~g19700)&(~g15257));
assign II32928 = ((~g24835));
assign g29016 = ((~g28672)&(~g13487));
assign g29314 = ((~II38471));
assign g27908 = (g13886&g27391);
assign g24758 = (g15618&g24111);
assign g13359 = ((~II20444));
assign II32697 = ((~g14280))|((~II32695));
assign II20467 = ((~g11263))|((~II20465));
assign II39635 = ((~g30055));
assign II21905 = ((~g13140));
assign g12305 = ((~g10593)&(~g10638)&(~g10670));
assign g8870 = ((~II16128));
assign g23837 = ((~II31071));
assign II32907 = ((~g24551));
assign g20188 = (g18593&g9425);
assign II24049 = ((~g16213));
assign II29903 = ((~g23134));
assign g30092 = (g29849&g11205);
assign II30901 = ((~g21974));
assign g22275 = ((~g20711));
assign g25590 = ((~II33415));
assign g13160 = ((~g8704)&(~g8717)&(~g8751));
assign g17145 = ((~g13971))|((~g13934));
assign II34244 = ((~g25253));
assign II39942 = ((~g30301));
assign g8491 = (g3566&g1618);
assign g16758 = ((~II22752));
assign g28167 = ((~g27456));
assign II39540 = ((~g29911))|((~II39539));
assign II33852 = ((~g25471));
assign g19231 = (g18363)|(g18441);
assign g26811 = ((~g15283)&(~g26279));
assign II29165 = ((~g20898));
assign g21747 = ((~g20228))|((~g6574));
assign g26631 = ((~g25746));
assign g22990 = ((~g21677)&(~g21078));
assign g13467 = ((~II20700));
assign II15654 = ((~g7085));
assign g30473 = (g30171&g11303);
assign g6079 = ((~II14584));
assign g29783 = ((~g29483)&(~g29235));
assign II16053 = ((~g6067));
assign g19575 = (g8194&g17307);
assign II28969 = ((~g21686));
assign g22267 = ((~g21731)&(~g20039));
assign II39821 = ((~g30267));
assign II14942 = ((~g2480));
assign II27074 = ((~g19238));
assign g15037 = ((~II21392));
assign g30826 = ((~II40730));
assign g12840 = ((~II19901));
assign g27336 = ((~g27088)&(~g26455));
assign II18311 = ((~g5668));
assign g18004 = ((~g14280));
assign g20941 = ((~g19724)&(~g17634));
assign g30792 = ((~II40634));
assign g10704 = (g3366&g5352);
assign g15869 = ((~g12657))|((~g6574));
assign g23111 = ((~g17091)&(~g21175));
assign g8498 = (g7085&g2309);
assign g30304 = ((~g13527)&(~g30007));
assign II37793 = ((~g28638));
assign II39005 = ((~g29507));
assign g11025 = ((~II17936));
assign g24351 = ((~II31727));
assign II25231 = ((~g18952));
assign g11535 = ((~II18581));
assign g15999 = ((~g12955))|((~g7230));
assign II31226 = ((~g22651));
assign II37056 = ((~g28082));
assign g28240 = ((~II36969));
assign g13191 = ((~g9484));
assign g24183 = ((~II31387));
assign II32333 = ((~g18131))|((~g23997));
assign g13107 = ((~g10822));
assign II16037 = ((~g6061));
assign g11726 = ((~g9676))|((~g3522));
assign II19883 = ((~g8550));
assign g26280 = ((~II34238));
assign g21528 = ((~II28061));
assign g18807 = ((~g15112));
assign g12409 = ((~II19557));
assign II23292 = ((~g13741));
assign g24435 = (g17151&g24168&g13649);
endmodule
