module s15850(
  blif_clk_net,
  blif_reset_net,
  g18,
  g27,
  g109,
  g741,
  g742,
  g743,
  g744,
  g872,
  g873,
  g877,
  g881,
  g1712,
  g1960,
  g1961,
  g2355,
  g2601,
  g2602,
  g2603,
  g2604,
  g2605,
  g2606,
  g2607,
  g2608,
  g2609,
  g2610,
  g2611,
  g2612,
  g2648,
  g2986,
  g3007,
  g3069,
  g4172,
  g4173,
  g4174,
  g4175,
  g4176,
  g4177,
  g4178,
  g4179,
  g4180,
  g4181,
  g4887,
  g4888,
  g5101,
  g5105,
  g5658,
  g5659,
  g5816,
  g6920,
  g6926,
  g6932,
  g6942,
  g6949,
  g6955,
  g7744,
  g8061,
  g8062,
  g8271,
  g8313,
  g8316,
  g8318,
  g8323,
  g8328,
  g8331,
  g8335,
  g8340,
  g8347,
  g8349,
  g8352,
  g8561,
  g8562,
  g8563,
  g8564,
  g8565,
  g8566,
  g8976,
  g8977,
  g8978,
  g8979,
  g8980,
  g8981,
  g8982,
  g8983,
  g8984,
  g8985,
  g8986,
  g9451,
  g9961,
  g10377,
  g10379,
  g10455,
  g10457,
  g10459,
  g10461,
  g10463,
  g10465,
  g10628,
  g10801,
  g11163,
  g11206,
  g11489);
input blif_clk_net;
input blif_reset_net;
input g18;
input g27;
input g109;
input g741;
input g742;
input g743;
input g744;
input g872;
input g873;
input g877;
input g881;
input g1712;
input g1960;
input g1961;
output g2355;
output g2601;
output g2602;
output g2603;
output g2604;
output g2605;
output g2606;
output g2607;
output g2608;
output g2609;
output g2610;
output g2611;
output g2612;
output g2648;
output g2986;
output g3007;
output g3069;
output g4172;
output g4173;
output g4174;
output g4175;
output g4176;
output g4177;
output g4178;
output g4179;
output g4180;
output g4181;
output g4887;
output g4888;
output g5101;
output g5105;
output g5658;
output g5659;
output g5816;
output g6920;
output g6926;
output g6932;
output g6942;
output g6949;
output g6955;
output g7744;
output g8061;
output g8062;
output g8271;
output g8313;
output g8316;
output g8318;
output g8323;
output g8328;
output g8331;
output g8335;
output g8340;
output g8347;
output g8349;
output g8352;
output g8561;
output g8562;
output g8563;
output g8564;
output g8565;
output g8566;
output g8976;
output g8977;
output g8978;
output g8979;
output g8980;
output g8981;
output g8982;
output g8983;
output g8984;
output g8985;
output g8986;
output g9451;
output g9961;
output g10377;
output g10379;
output g10455;
output g10457;
output g10459;
output g10461;
output g10463;
output g10465;
output g10628;
output g10801;
output g11163;
output g11206;
output g11489;
reg g30;
reg g31;
reg g32;
reg g33;
reg g34;
reg g35;
reg g36;
reg g37;
reg g38;
reg g39;
reg g40;
reg g41;
reg g42;
reg g43;
reg g44;
reg g45;
reg g46;
reg g47;
reg g48;
reg g82;
reg g83;
reg g84;
reg g85;
reg g86;
reg g87;
reg g88;
reg g89;
reg g90;
reg g91;
reg g92;
reg g93;
reg g94;
reg g95;
reg g96;
reg g99;
reg g100;
reg g101;
reg g102;
reg g103;
reg g104;
reg g28;
reg g29;
reg g898;
reg g901;
reg g904;
reg g907;
reg g910;
reg g913;
reg g916;
reg g919;
reg g922;
reg g925;
reg g971;
reg g976;
reg g981;
reg g986;
reg g944;
reg g947;
reg g950;
reg g953;
reg g956;
reg g959;
reg g962;
reg g965;
reg g968;
reg g886;
reg g889;
reg g892;
reg g895;
reg g928;
reg g932;
reg g936;
reg g940;
reg g883;
reg g882;
reg g878;
reg g876;
reg g757;
reg g755;
reg g756;
reg g745;
reg g746;
reg g750;
reg g754;
reg g758;
reg g762;
reg g766;
reg g770;
reg g774;
reg g778;
reg g782;
reg g786;
reg g790;
reg g865;
reg g794;
reg g798;
reg g802;
reg g806;
reg g810;
reg g814;
reg g818;
reg g822;
reg g826;
reg g829;
reg g833;
reg g837;
reg g841;
reg g845;
reg g849;
reg g853;
reg g857;
reg g861;
reg g874;
reg g868;
reg g875;
reg g869;
reg g590;
reg g584;
reg g585;
reg g586;
reg g587;
reg g588;
reg g589;
reg g578;
reg g579;
reg g580;
reg g581;
reg g582;
reg g583;
reg g253;
reg g256;
reg g257;
reg g258;
reg g259;
reg g260;
reg g261;
reg g262;
reg g254;
reg g255;
reg g143;
reg g166;
reg g139;
reg g135;
reg g131;
reg g127;
reg g170;
reg g174;
reg g162;
reg g158;
reg g153;
reg g148;
reg g178;
reg g182;
reg g126;
reg g263;
reg g266;
reg g269;
reg g272;
reg g275;
reg g278;
reg g281;
reg g284;
reg g287;
reg g290;
reg g293;
reg g296;
reg g299;
reg g302;
reg g123;
reg g119;
reg g611;
reg g617;
reg g591;
reg g599;
reg g605;
reg g630;
reg g631;
reg g632;
reg g635;
reg g627;
reg g636;
reg g639;
reg g622;
reg g643;
reg g646;
reg g650;
reg g654;
reg g658;
reg g668;
reg g677;
reg g686;
reg g695;
reg g704;
reg g713;
reg g722;
reg g731;
reg g664;
reg g673;
reg g682;
reg g691;
reg g700;
reg g709;
reg g718;
reg g727;
reg g736;
reg g8;
reg g17;
reg g481;
reg g486;
reg g491;
reg g496;
reg g501;
reg g506;
reg g511;
reg g516;
reg g476;
reg g542;
reg g538;
reg g534;
reg g530;
reg g525;
reg g521;
reg g456;
reg g461;
reg g466;
reg g471;
reg g305;
reg g315;
reg g318;
reg g321;
reg g324;
reg g327;
reg g330;
reg g333;
reg g309;
reg g312;
reg g426;
reg g386;
reg g391;
reg g396;
reg g401;
reg g406;
reg g411;
reg g416;
reg g421;
reg g452;
reg g448;
reg g444;
reg g440;
reg g435;
reg g431;
reg g369;
reg g374;
reg g378;
reg g382;
reg g336;
reg g348;
reg g351;
reg g354;
reg g357;
reg g360;
reg g363;
reg g366;
reg g342;
reg g339;
reg g345;
reg g49;
reg g52;
reg g55;
reg g58;
reg g61;
reg g64;
reg g67;
reg g70;
reg g73;
reg g76;
reg g79;
reg g113;
reg g114;
reg g1955;
reg g1956;
reg g1957;
reg g1700;
reg g1696;
reg g1703;
reg g1710;
reg g1713;
reg g1718;
reg g1766;
reg g1771;
reg g1776;
reg g1781;
reg g1786;
reg g1791;
reg g1796;
reg g1801;
reg g1806;
reg g1711;
reg g1834;
reg g1840;
reg g1814;
reg g1822;
reg g1828;
reg g1848;
reg g1849;
reg g1850;
reg g1853;
reg g1845;
reg g1854;
reg g1857;
reg g1861;
reg g1864;
reg g1868;
reg g1872;
reg g1882;
reg g1891;
reg g1900;
reg g1909;
reg g1918;
reg g1927;
reg g1936;
reg g1945;
reg g1878;
reg g1887;
reg g1896;
reg g1905;
reg g1914;
reg g1923;
reg g1932;
reg g1941;
reg g1950;
reg g16;
reg g7;
reg g1736;
reg g1737;
reg g1648;
reg g1651;
reg g1642;
reg g1645;
reg g1610;
reg g1765;
reg g1811;
reg g1721;
reg g1724;
reg g1727;
reg g1730;
reg g1733;
reg g1738;
reg g1741;
reg g1744;
reg g1747;
reg g1750;
reg g1753;
reg g1756;
reg g1759;
reg g1762;
reg g1958;
reg g1810;
reg g1959;
reg g1707;
reg g1690;
reg g1170;
reg g1173;
reg g1176;
reg g1179;
reg g1182;
reg g1185;
reg g1188;
reg g1191;
reg g1194;
reg g1197;
reg g1200;
reg g1203;
reg g1169;
reg g108;
reg g1336;
reg g1341;
reg g1346;
reg g1351;
reg g1206;
reg g1361;
reg g1360;
reg g1216;
reg g1217;
reg g1212;
reg g1209;
reg g1215;
reg g1357;
reg g1289;
reg g1275;
reg g1235;
reg g1240;
reg g1245;
reg g1250;
reg g1255;
reg g1260;
reg g1265;
reg g1270;
reg g1304;
reg g1300;
reg g1296;
reg g1292;
reg g1284;
reg g1280;
reg g1218;
reg g1223;
reg g1227;
reg g1231;
reg g1356;
reg g1317;
reg g1314;
reg g1318;
reg g1321;
reg g1324;
reg g1327;
reg g1330;
reg g1333;
reg g1308;
reg g1311;
reg g1035;
reg g1047;
reg g1050;
reg g1053;
reg g1056;
reg g1059;
reg g1062;
reg g1065;
reg g1038;
reg g1041;
reg g1044;
reg g1068;
reg g1080;
reg g1083;
reg g1086;
reg g1089;
reg g1092;
reg g1095;
reg g1098;
reg g1074;
reg g1071;
reg g1077;
reg g1027;
reg g995;
reg g991;
reg g1003;
reg g999;
reg g1011;
reg g1007;
reg g1019;
reg g1015;
reg g1023;
reg g1032;
reg g105;
reg g1117;
reg g1121;
reg g1125;
reg g1129;
reg g1133;
reg g1137;
reg g1141;
reg g1145;
reg g1113;
reg g1166;
reg g1163;
reg g1160;
reg g1157;
reg g1153;
reg g1149;
reg g1101;
reg g1104;
reg g1107;
reg g1110;
reg g1618;
reg g1615;
reg g1621;
reg g1624;
reg g1627;
reg g1630;
reg g1633;
reg g1636;
reg g1639;
reg g1512;
reg g1448;
reg g1444;
reg g1440;
reg g1436;
reg g1432;
reg g1403;
reg g1428;
reg g1407;
reg g1424;
reg g1411;
reg g1419;
reg g1515;
reg g1520;
reg g1415;
reg g1453;
reg g1458;
reg g1462;
reg g1466;
reg g1470;
reg g1474;
reg g1478;
reg g1482;
reg g1486;
reg g1490;
reg g1494;
reg g1499;
reg g1504;
reg g1508;
reg g1393;
reg g1394;
reg g115;
reg g201;
reg g1374;
reg g197;
reg g1389;
reg g192;
reg g1397;
reg g248;
reg g1400;
reg g243;
reg g1362;
reg g237;
reg g1365;
reg g231;
reg g1368;
reg g225;
reg g1371;
reg g219;
reg g1377;
reg g213;
reg g1380;
reg g207;
reg g1383;
reg g186;
reg g1386;
reg g4;
reg g12;
reg g1;
reg g9;
reg g1527;
reg g1524;
reg g1528;
reg g1531;
reg g1534;
reg g1537;
reg g1540;
reg g1543;
reg g1546;
reg g1549;
reg g1552;
reg g1555;
reg g1558;
reg g1561;
reg g1564;
reg g1570;
reg g1567;
reg g1571;
reg g1574;
reg g1577;
reg g1580;
reg g1583;
reg g1586;
reg g1589;
reg g1592;
reg g1595;
reg g1598;
reg g1601;
reg g1604;
reg g1607;
reg g1654;
reg g1657;
reg g1660;
reg g1663;
reg g1666;
reg g1669;
reg g1672;
reg g1675;
reg g1678;
reg g1681;
reg g1684;
reg g1687;
reg g546;
reg g554;
reg g557;
reg g560;
reg g563;
reg g566;
reg g569;
reg g572;
reg g575;
reg g549;
reg g552;
reg g553;
reg g23;
reg g26;
wire g2171;
wire g3491;
wire g2000;
wire g10722;
wire II12647;
wire g6579;
wire g10241;
wire II13463;
wire II10924;
wire II12216;
wire II14835;
wire g10306;
wire g10861;
wire g4866;
wire g8600;
wire g3783;
wire g8117;
wire g8508;
wire g8487;
wire g6136;
wire g10300;
wire II4783;
wire g7555;
wire g8588;
wire g11145;
wire g7570;
wire g7881;
wire g7658;
wire g2776;
wire II12226;
wire g9834;
wire g9621;
wire g6426;
wire g8278;
wire II10349;
wire II8711;
wire II7405;
wire g8946;
wire g9700;
wire g10764;
wire II5315;
wire g8932;
wire II7562;
wire g4960;
wire g9338;
wire g6045;
wire g3221;
wire II5891;
wire g10695;
wire g7246;
wire g2039;
wire II7432;
wire g11192;
wire II16051;
wire g5845;
wire g2321;
wire II5095;
wire II10228;
wire g7440;
wire II5689;
wire g2662;
wire g7600;
wire II15871;
wire g8801;
wire g7756;
wire g5119;
wire g5099;
wire g7636;
wire II7441;
wire g10310;
wire g4097;
wire II10039;
wire g5778;
wire g8641;
wire g9606;
wire II16847;
wire g10947;
wire g4157;
wire g8938;
wire g5913;
wire g9901;
wire g6544;
wire g5589;
wire g10743;
wire gbuf10;
wire II11907;
wire g4276;
wire g10950;
wire g2651;
wire g8941;
wire g7521;
wire g6358;
wire g10560;
wire g4897;
wire g3638;
wire II15542;
wire II11440;
wire II16332;
wire g9830;
wire g11259;
wire g10668;
wire g9717;
wire II16161;
wire g8717;
wire g10877;
wire g6890;
wire g10732;
wire g9809;
wire gbuf3;
wire II8562;
wire g11545;
wire g10872;
wire II17407;
wire g10783;
wire II6631;
wire g2503;
wire g8106;
wire II7109;
wire g2135;
wire g10230;
wire II15187;
wire II5192;
wire g6114;
wire II9804;
wire g11232;
wire II16550;
wire g6847;
wire g6818;
wire g10495;
wire g10685;
wire g5491;
wire g10882;
wire g8645;
wire II11436;
wire g10186;
wire g4883;
wire II17730;
wire g6015;
wire g7136;
wire g4939;
wire g5726;
wire g2177;
wire II16407;
wire II15281;
wire g9962;
wire g8885;
wire g6827;
wire g8143;
wire g10778;
wire g5673;
wire g11650;
wire g8130;
wire II10507;
wire g5295;
wire g6743;
wire g6101;
wire II6543;
wire II8256;
wire g11472;
wire g8123;
wire g7569;
wire g3748;
wire g6279;
wire g9109;
wire II12678;
wire g7942;
wire g5318;
wire II11427;
wire g4919;
wire II11417;
wire g6594;
wire g8817;
wire II16540;
wire g8032;
wire II17243;
wire g9738;
wire g6155;
wire g11584;
wire g7914;
wire g5602;
wire g1976;
wire II4941;
wire g9665;
wire g8704;
wire II9647;
wire II13544;
wire g2087;
wire II15539;
wire II11773;
wire g6333;
wire II13858;
wire g2315;
wire g6108;
wire II8982;
wire g6389;
wire g10270;
wire g4899;
wire g7264;
wire II12406;
wire g3385;
wire g6364;
wire g8219;
wire g11575;
wire g3200;
wire g5185;
wire g4459;
wire g9347;
wire g4717;
wire g8384;
wire g10217;
wire II15314;
wire g10025;
wire g4413;
wire g4127;
wire g10117;
wire g8804;
wire g5947;
wire II9259;
wire II5485;
wire II13933;
wire g1982;
wire II5391;
wire g10125;
wire II9893;
wire g7818;
wire g5935;
wire g10134;
wire g6086;
wire g7297;
wire g11266;
wire g11331;
wire g5258;
wire II5500;
wire g2941;
wire g3990;
wire g2727;
wire g10894;
wire g2340;
wire g2054;
wire g7132;
wire II16766;
wire g7797;
wire II13714;
wire g1989;
wire g9709;
wire g9360;
wire g8210;
wire g6822;
wire II8831;
wire g7409;
wire g10400;
wire II15060;
wire g8044;
wire II5792;
wire II7665;
wire II6901;
wire g11284;
wire g2984;
wire II14449;
wire g8137;
wire g5512;
wire g10405;
wire g4461;
wire g4168;
wire g6488;
wire II14271;
wire g4720;
wire g7588;
wire g6150;
wire II6643;
wire g7537;
wire g9868;
wire g6662;
wire g5489;
wire g6269;
wire g3109;
wire g9582;
wire g2181;
wire g4999;
wire g11032;
wire II8333;
wire g7962;
wire g2328;
wire g9696;
wire g5305;
wire II9341;
wire g9357;
wire II7303;
wire II13962;
wire II13341;
wire g9914;
wire g8461;
wire g2157;
wire II17337;
wire g2014;
wire g11633;
wire II12085;
wire g6536;
wire g9271;
wire g11169;
wire g8556;
wire g10201;
wire g4064;
wire g8250;
wire g3807;
wire g10453;
wire II14506;
wire g6900;
wire g2669;
wire g5074;
wire II5085;
wire g3213;
wire II5459;
wire II10042;
wire g9683;
wire g11344;
wire g7681;
wire g2733;
wire II11330;
wire II14855;
wire II6861;
wire II9279;
wire g2462;
wire II17563;
wire g2246;
wire g11506;
wire g11484;
wire g4777;
wire II6414;
wire II9992;
wire II7577;
wire g5525;
wire g6654;
wire g11006;
wire g10328;
wire g5815;
wire g3991;
wire II15858;
wire g4637;
wire g7364;
wire g2025;
wire II10048;
wire g11613;
wire II13430;
wire g9825;
wire II7487;
wire g4285;
wire II11524;
wire g7316;
wire g5274;
wire g2614;
wire II15042;
wire g6961;
wire g10527;
wire g7339;
wire g2211;
wire g5210;
wire g11045;
wire g8206;
wire g6225;
wire g3051;
wire II9680;
wire g5820;
wire II16203;
wire g7747;
wire g10279;
wire g4468;
wire g3066;
wire II6225;
wire g5268;
wire g6416;
wire g5038;
wire g8159;
wire g3463;
wire g7896;
wire II16360;
wire II14315;
wire g4508;
wire g11342;
wire II10801;
wire g7386;
wire g10373;
wire g8293;
wire II15778;
wire g7449;
wire II5237;
wire II15311;
wire II12193;
wire g7024;
wire II16979;
wire g10969;
wire II9639;
wire g6176;
wire II9020;
wire g4972;
wire II10398;
wire II13523;
wire II10834;
wire g6909;
wire g11081;
wire II5064;
wire g2683;
wire II5667;
wire g10762;
wire g11080;
wire II6742;
wire g3398;
wire g7787;
wire g4267;
wire II11034;
wire g3144;
wire II5510;
wire g10972;
wire II13230;
wire g7143;
wire g10332;
wire II12550;
wire g10770;
wire g6884;
wire II16679;
wire II15962;
wire g3475;
wire g11491;
wire g7147;
wire g6049;
wire II15861;
wire g10007;
wire II6156;
wire II7877;
wire g7593;
wire g11550;
wire g9111;
wire g7676;
wire g4732;
wire II15256;
wire g10854;
wire II13738;
wire g10333;
wire II11992;
wire g5894;
wire II17453;
wire g10384;
wire g2334;
wire g11260;
wire II13695;
wire g10616;
wire II10958;
wire g2990;
wire g3697;
wire II10546;
wire g10543;
wire g7734;
wire II17225;
wire II6031;
wire II10598;
wire g7761;
wire g6252;
wire II13831;
wire g4435;
wire II10421;
wire g8891;
wire II5441;
wire g5766;
wire II13083;
wire g4283;
wire g10165;
wire II9240;
wire g4824;
wire g7075;
wire g2864;
wire II10168;
wire g10545;
wire g7049;
wire g11108;
wire g8640;
wire g6569;
wire g9919;
wire g5624;
wire g2771;
wire g8844;
wire g8837;
wire g8664;
wire g7137;
wire II9550;
wire g2482;
wire II6454;
wire g11022;
wire g11224;
wire g7390;
wire II5662;
wire g4219;
wire g4790;
wire g9876;
wire II13125;
wire g3517;
wire II15088;
wire II11397;
wire g9448;
wire II11149;
wire II15782;
wire g3585;
wire II16708;
wire g7307;
wire g10140;
wire g11324;
wire II5373;
wire g4170;
wire II5632;
wire g6804;
wire g10729;
wire g2253;
wire g7908;
wire g3375;
wire II11176;
wire g3874;
wire g11196;
wire II6598;
wire II8671;
wire II15403;
wire II9352;
wire g6899;
wire g10750;
wire II9938;
wire g10692;
wire g5010;
wire g5650;
wire II10816;
wire g6670;
wire g6465;
wire II17149;
wire g5251;
wire g10092;
wire g10043;
wire g5405;
wire II10090;
wire g10503;
wire g4678;
wire g5630;
wire g7709;
wire g3631;
wire g3726;
wire g7950;
wire II5403;
wire II12613;
wire II16239;
wire II15085;
wire g11295;
wire II12478;
wire g6260;
wire II13272;
wire II7288;
wire g6679;
wire II14094;
wire g2373;
wire II17461;
wire g6064;
wire g2918;
wire g2959;
wire II16613;
wire g4873;
wire II14228;
wire g7330;
wire g3945;
wire g4596;
wire g4613;
wire g11616;
wire g6771;
wire g11241;
wire g8131;
wire g7610;
wire g10265;
wire g8446;
wire g8781;
wire g9426;
wire g6553;
wire g10794;
wire II13239;
wire II8869;
wire g4048;
wire II14522;
wire g8426;
wire II14263;
wire II12989;
wire II8154;
wire g11304;
wire g5882;
wire g4840;
wire g5486;
wire II11058;
wire II6085;
wire II8303;
wire g2647;
wire II11228;
wire II13723;
wire g8152;
wire II8178;
wire g3118;
wire g9566;
wire II9559;
wire g8501;
wire g3721;
wire g2406;
wire g5747;
wire g7268;
wire II6996;
wire g9366;
wire g6308;
wire g7656;
wire g11230;
wire g8434;
wire II12832;
wire g2203;
wire II7701;
wire II8320;
wire II8240;
wire g2541;
wire II6488;
wire g1998;
wire g3228;
wire g3903;
wire g2354;
wire g5864;
wire II10702;
wire II8631;
wire g8962;
wire II16095;
wire II15729;
wire g7070;
wire g3076;
wire II5135;
wire II6406;
wire g7894;
wire II16629;
wire g5395;
wire II13589;
wire II8436;
wire g5689;
wire g7191;
wire g9716;
wire g11046;
wire II12535;
wire g2832;
wire II7354;
wire II13669;
wire II7633;
wire II17513;
wire II8590;
wire II13822;
wire II11106;
wire g4054;
wire II12143;
wire g2964;
wire g10348;
wire II10666;
wire g10177;
wire g11586;
wire g10575;
wire II9199;
wire g7213;
wire g10175;
wire g8768;
wire g5984;
wire g7358;
wire g6094;
wire II5015;
wire g9124;
wire g9262;
wire g4213;
wire g6924;
wire II7779;
wire g6070;
wire g11222;
wire g4730;
wire g3459;
wire g3291;
wire II9008;
wire g9595;
wire g7603;
wire g4094;
wire g7884;
wire II12127;
wire II8513;
wire II14236;
wire g6541;
wire II5588;
wire g6995;
wire g3435;
wire II12916;
wire II13096;
wire g10880;
wire g5693;
wire g2222;
wire g11311;
wire II6439;
wire g2891;
wire g7972;
wire g10204;
wire g2369;
wire g7011;
wire g6970;
wire II5943;
wire II11713;
wire g8418;
wire II4906;
wire g10667;
wire II5989;
wire II11980;
wire g6248;
wire g4307;
wire g8883;
wire g10440;
wire g10507;
wire g4343;
wire II16802;
wire II13391;
wire II9001;
wire g11237;
wire g8362;
wire g5875;
wire g10194;
wire g10536;
wire g11248;
wire g11070;
wire II14613;
wire g7926;
wire II12773;
wire g5514;
wire g8069;
wire g11557;
wire g7227;
wire g9512;
wire g2274;
wire II6178;
wire II12239;
wire II9162;
wire II17185;
wire g2548;
wire g11306;
wire g11062;
wire g5026;
wire g5682;
wire II11405;
wire g4395;
wire g8187;
wire g3685;
wire II15356;
wire g8846;
wire g2213;
wire II5734;
wire g5547;
wire II12770;
wire g10339;
wire II8449;
wire II6958;
wire g3343;
wire II6528;
wire II10633;
wire g11155;
wire II9302;
wire g5446;
wire g6309;
wire g9758;
wire g10902;
wire g11033;
wire g3068;
wire g10466;
wire g7377;
wire g2858;
wire g9029;
wire g7791;
wire g6395;
wire II15412;
wire g4115;
wire g10188;
wire II17402;
wire g7531;
wire g3332;
wire g3396;
wire II11315;
wire g5477;
wire g3095;
wire g10365;
wire g5062;
wire g3437;
wire g10624;
wire g8788;
wire g11630;
wire II10563;
wire g7185;
wire g5149;
wire g7538;
wire II5231;
wire g5540;
wire g5888;
wire g3911;
wire II11132;
wire g3760;
wire g4321;
wire g2239;
wire g6186;
wire g11363;
wire g5277;
wire II13571;
wire g3767;
wire II12583;
wire g8727;
wire II11786;
wire g8557;
wire g7022;
wire II7790;
wire g5197;
wire g5217;
wire g2111;
wire II10736;
wire g7935;
wire g4601;
wire g6200;
wire g3792;
wire g3383;
wire II6167;
wire g8402;
wire g7678;
wire g10594;
wire g9751;
wire II12020;
wire II9795;
wire g9385;
wire II17504;
wire g4669;
wire II10519;
wire g9936;
wire g3429;
wire g7458;
wire g6588;
wire g2079;
wire II5080;
wire II12652;
wire g3327;
wire II17307;
wire II9872;
wire g7810;
wire II6825;
wire II7225;
wire II14439;
wire g7056;
wire g4221;
wire II16510;
wire g10911;
wire g6524;
wire II5120;
wire g6196;
wire II9869;
wire II6894;
wire g10581;
wire g6941;
wire g6077;
wire II16871;
wire g9052;
wire II4891;
wire g11455;
wire g9667;
wire g6685;
wire g9956;
wire g9766;
wire II10308;
wire g3405;
wire g2306;
wire g8072;
wire g6392;
wire II15127;
wire g10438;
wire g5231;
wire II15275;
wire II7393;
wire g4309;
wire g2509;
wire g5995;
wire II6971;
wire g5782;
wire II9786;
wire II14087;
wire g10599;
wire g8550;
wire g10475;
wire g4237;
wire g7937;
wire II6061;
wire II12809;
wire g2571;
wire II17662;
wire g3626;
wire II5646;
wire g9257;
wire g6530;
wire II6124;
wire g8953;
wire II8651;
wire g5069;
wire g2456;
wire II7360;
wire g4226;
wire g8926;
wire II16277;
wire II12786;
wire II11674;
wire II6118;
wire II9232;
wire g2043;
wire II12526;
wire g4411;
wire g4755;
wire II8311;
wire g10699;
wire g9533;
wire g6322;
wire g10935;
wire g6207;
wire g9598;
wire g11013;
wire II14884;
wire II17543;
wire II13406;
wire g3415;
wire II7863;
wire g8163;
wire g10019;
wire II15389;
wire g7702;
wire g3120;
wire II10021;
wire g8167;
wire II16220;
wire II13682;
wire g2554;
wire g8341;
wire g6698;
wire g11377;
wire II6385;
wire g10515;
wire g7752;
wire g10483;
wire II16331;
wire g9742;
wire II6025;
wire g10427;
wire g4196;
wire g10649;
wire II9126;
wire g4457;
wire g11167;
wire g9351;
wire II9754;
wire g5574;
wire II11596;
wire g11388;
wire II6665;
wire II10678;
wire g10806;
wire g5202;
wire g10524;
wire g7201;
wire g11400;
wire II12508;
wire g6799;
wire g10255;
wire g5526;
wire g6435;
wire g11431;
wire II12344;
wire II9915;
wire g7906;
wire g7544;
wire g8710;
wire II11112;
wire g10396;
wire II5652;
wire g8081;
wire II16058;
wire II10015;
wire g10727;
wire II13869;
wire g4513;
wire g2411;
wire g11515;
wire g7726;
wire II6467;
wire g9643;
wire g6858;
wire g11316;
wire g6302;
wire g8052;
wire g8005;
wire g4388;
wire g4312;
wire g6706;
wire II11238;
wire g11051;
wire g9950;
wire g10287;
wire II17198;
wire II10120;
wire g10321;
wire II6173;
wire g11651;
wire II7163;
wire g10679;
wire II16190;
wire g8354;
wire II7964;
wire g5178;
wire II17340;
wire g5125;
wire II8136;
wire II17282;
wire g11188;
wire g4206;
wire g9525;
wire II10003;
wire II8763;
wire g7320;
wire g9659;
wire g4997;
wire g4161;
wire g5228;
wire g6660;
wire g2260;
wire II9816;
wire g10229;
wire g11541;
wire g6472;
wire II9576;
wire g6764;
wire II12466;
wire g6747;
wire g2379;
wire g5537;
wire II8414;
wire g3044;
wire g6314;
wire II17152;
wire g10630;
wire g9672;
wire g6368;
wire g2475;
wire II8544;
wire II6209;
wire g3262;
wire II11841;
wire g5120;
wire II11024;
wire g4482;
wire II17176;
wire g4948;
wire g4901;
wire g11621;
wire g4764;
wire g4559;
wire g7053;
wire g8327;
wire g4067;
wire g10739;
wire g8994;
wire II9498;
wire II13840;
wire II16775;
wire g11102;
wire g10308;
wire g10512;
wire g10675;
wire g4503;
wire II12463;
wire II10129;
wire g10294;
wire II7825;
wire II11737;
wire II5789;
wire II5171;
wire gbuf5;
wire g6841;
wire g7066;
wire g9100;
wire g5003;
wire g6871;
wire II11858;
wire II10384;
wire II13078;
wire g3817;
wire g5804;
wire g6617;
wire g10447;
wire II15989;
wire g5787;
wire II6277;
wire g10639;
wire g7803;
wire g9894;
wire II5979;
wire II7402;
wire g9776;
wire II17531;
wire II11286;
wire g10926;
wire g4095;
wire II15359;
wire II10132;
wire g6736;
wire g10301;
wire II15365;
wire g4240;
wire g2083;
wire g8288;
wire g3257;
wire g8471;
wire g2907;
wire g6255;
wire g9316;
wire g11438;
wire II6793;
wire g6792;
wire g9421;
wire II17324;
wire II8796;
wire g11207;
wire g5170;
wire g10730;
wire II11563;
wire g10825;
wire g9602;
wire g6217;
wire g11336;
wire g11069;
wire g5847;
wire II6826;
wire g9873;
wire II15759;
wire g2819;
wire g8413;
wire g8065;
wire II12634;
wire II8677;
wire II9391;
wire g6227;
wire II5539;
wire g9449;
wire g6838;
wire II10198;
wire II14330;
wire II8495;
wire II6052;
wire g3507;
wire g8526;
wire g10350;
wire g10159;
wire g5209;
wire II8788;
wire g2342;
wire II7131;
wire g9267;
wire g9848;
wire g2749;
wire II12415;
wire g6162;
wire g2523;
wire g8247;
wire g9925;
wire g8638;
wire II7837;
wire g10870;
wire II7899;
wire g3252;
wire II5105;
wire g8375;
wire g5763;
wire II10237;
wire g5041;
wire II8085;
wire g11059;
wire II14382;
wire g8877;
wire g4804;
wire g5281;
wire g2164;
wire g8301;
wire g9650;
wire g4545;
wire g6000;
wire g2125;
wire g11485;
wire g7997;
wire g6628;
wire g4564;
wire g5424;
wire II5414;
wire g4056;
wire g10420;
wire g2115;
wire II15497;
wire II7984;
wire g6739;
wire g11216;
wire II16172;
wire g4328;
wire g4606;
wire II7938;
wire g3828;
wire II4951;
wire g11274;
wire g6112;
wire II11214;
wire II6832;
wire II10069;
wire II5204;
wire g10472;
wire g3773;
wire g4332;
wire g9722;
wire g10378;
wire II11743;
wire II13379;
wire g7107;
wire g6099;
wire II15362;
wire g6362;
wire g5051;
wire II16209;
wire g8382;
wire II9531;
wire g5183;
wire g4715;
wire II8576;
wire II15880;
wire g7500;
wire g7928;
wire g6140;
wire g3757;
wire II15974;
wire II15220;
wire g9355;
wire II12060;
wire g10697;
wire II5006;
wire g9027;
wire g5987;
wire II9984;
wire g2586;
wire g9274;
wire II13335;
wire II8247;
wire g7236;
wire g7295;
wire g3718;
wire g9987;
wire g6157;
wire g6335;
wire g3804;
wire II7311;
wire g8702;
wire II13766;
wire g10547;
wire g6294;
wire g4062;
wire g6250;
wire g7795;
wire g11573;
wire g11501;
wire g10493;
wire II16376;
wire g4129;
wire g8815;
wire g11161;
wire g8653;
wire II5982;
wire II5336;
wire g4116;
wire g8436;
wire II17568;
wire II10557;
wire g9707;
wire II7833;
wire g6050;
wire g8108;
wire g6745;
wire g7326;
wire g11268;
wire g7707;
wire g11039;
wire II10931;
wire g5151;
wire II15980;
wire g2943;
wire g11655;
wire g9963;
wire g8018;
wire g3728;
wire g5982;
wire g4786;
wire II13595;
wire g8944;
wire g2089;
wire II5502;
wire g8698;
wire g5028;
wire II11620;
wire g9862;
wire g5443;
wire II8481;
wire II5801;
wire II10391;
wire g7021;
wire II9077;
wire g6731;
wire II13267;
wire g9584;
wire II13357;
wire g6406;
wire g5147;
wire g9916;
wire g6298;
wire II6648;
wire g5552;
wire II6010;
wire II12574;
wire II11635;
wire g8735;
wire II13729;
wire g3206;
wire g2744;
wire II6381;
wire g2913;
wire g8054;
wire g2167;
wire g7535;
wire II9099;
wire II16944;
wire II11088;
wire II8739;
wire II6867;
wire g5949;
wire II12580;
wire II6531;
wire II7070;
wire g11600;
wire g3107;
wire g4722;
wire g4967;
wire g5668;
wire II14373;
wire g8281;
wire g6593;
wire g7960;
wire II16111;
wire II6784;
wire II7426;
wire g2230;
wire II15669;
wire II9144;
wire g11018;
wire g9727;
wire g6259;
wire g10160;
wire g7985;
wire II11611;
wire II16045;
wire II16543;
wire g5288;
wire II17761;
wire g8149;
wire g7711;
wire g6340;
wire II17052;
wire g10402;
wire II11272;
wire g10269;
wire II11162;
wire g10260;
wire g8603;
wire g5791;
wire II6217;
wire II12790;
wire g11263;
wire II9424;
wire g8171;
wire g9364;
wire g4608;
wire g5632;
wire g7586;
wire g4560;
wire g3209;
wire II4943;
wire g9858;
wire g10470;
wire g11631;
wire II17482;
wire g8709;
wire g2072;
wire g9311;
wire g6902;
wire g10661;
wire II11204;
wire g6263;
wire g8197;
wire g5706;
wire II9632;
wire g8652;
wire II7719;
wire g7777;
wire II15452;
wire g10570;
wire g4933;
wire II6350;
wire g10258;
wire g8485;
wire g8647;
wire g10319;
wire g7878;
wire g2632;
wire g9536;
wire II16691;
wire g7549;
wire g9818;
wire g9836;
wire g6351;
wire II6535;
wire II12901;
wire g11200;
wire II11293;
wire g7442;
wire g7754;
wire g6074;
wire II8805;
wire g7113;
wire g5519;
wire g3862;
wire II16181;
wire g9839;
wire g10754;
wire g2160;
wire II13612;
wire II15461;
wire g7634;
wire g4162;
wire g2002;
wire g4871;
wire g8936;
wire g2989;
wire g5227;
wire g7848;
wire g4506;
wire II16008;
wire g8643;
wire g10058;
wire g7883;
wire II16193;
wire g8488;
wire II10331;
wire g3393;
wire g11060;
wire g3368;
wire g10949;
wire g5915;
wire g9623;
wire g10741;
wire g2106;
wire g6032;
wire g9309;
wire II11489;
wire g2155;
wire g8141;
wire II14361;
wire g9832;
wire g11462;
wire g11199;
wire g4549;
wire g4524;
wire g4274;
wire g5117;
wire g2244;
wire g11029;
wire II10150;
wire II6207;
wire II4938;
wire II12069;
wire g8753;
wire II10538;
wire g10232;
wire II11689;
wire g10154;
wire II5528;
wire II6549;
wire g3703;
wire II6137;
wire II12481;
wire g9903;
wire g10247;
wire g5655;
wire II9317;
wire g10326;
wire g8315;
wire g8001;
wire g2653;
wire g10316;
wire g8959;
wire II10317;
wire g11234;
wire g11239;
wire g7616;
wire g8518;
wire g4478;
wire g9706;
wire g4989;
wire g6796;
wire g2956;
wire II8337;
wire g4385;
wire g8011;
wire g2418;
wire II9177;
wire g4210;
wire g6276;
wire g4372;
wire II4924;
wire g3742;
wire g3538;
wire g6475;
wire g6118;
wire g6829;
wire II5970;
wire g8121;
wire g5675;
wire II12019;
wire g9611;
wire g5530;
wire g6124;
wire g6382;
wire g5774;
wire II15054;
wire g11256;
wire g4553;
wire g2774;
wire g10879;
wire g2175;
wire g7244;
wire g6741;
wire II11519;
wire g11190;
wire II6982;
wire g2881;
wire g11470;
wire II16853;
wire g3633;
wire g6931;
wire g11297;
wire II15200;
wire g3733;
wire II6448;
wire g4428;
wire g2758;
wire g9223;
wire g10505;
wire II6391;
wire II14979;
wire g2645;
wire g10760;
wire II6347;
wire II12115;
wire g10737;
wire g5012;
wire II17764;
wire g2124;
wire g3876;
wire g7745;
wire g5256;
wire II5421;
wire g8133;
wire II16670;
wire II16108;
wire g8806;
wire II12205;
wire g10792;
wire g9874;
wire g3735;
wire g2971;
wire g8720;
wire g6199;
wire II8614;
wire II6183;
wire II13545;
wire g6704;
wire g4914;
wire II13457;
wire II6240;
wire II17365;
wire II7760;
wire II6188;
wire g6133;
wire II12046;
wire II5240;
wire g8400;
wire g9489;
wire g11194;
wire II8865;
wire II15215;
wire II6247;
wire g4681;
wire g6439;
wire g9345;
wire g6213;
wire g11326;
wire g8024;
wire g9846;
wire g4819;
wire g3142;
wire II6398;
wire g2826;
wire II7680;
wire II7064;
wire g6844;
wire g6893;
wire g11290;
wire g10857;
wire g9572;
wire II7244;
wire g11411;
wire II14080;
wire II15491;
wire g5745;
wire II5031;
wire II13791;
wire II14265;
wire g11105;
wire g3513;
wire g7305;
wire g11414;
wire g2939;
wire g8967;
wire g7512;
wire g8631;
wire II17687;
wire g6057;
wire g6571;
wire g2208;
wire g6447;
wire g8511;
wire II11043;
wire g2045;
wire g7110;
wire g5637;
wire g2916;
wire g1969;
wire g3751;
wire g10501;
wire II7556;
wire II5952;
wire II5450;
wire g4471;
wire g10115;
wire g2446;
wire g10937;
wire g7947;
wire II15672;
wire g8310;
wire g7453;
wire g8795;
wire g8960;
wire g10720;
wire g8338;
wire g5880;
wire g10863;
wire g3905;
wire II7973;
wire g8333;
wire II12354;
wire g9927;
wire g8623;
wire g5308;
wire g8276;
wire g8295;
wire g6824;
wire g4353;
wire II6944;
wire g2544;
wire g6870;
wire II7752;
wire II4996;
wire g11067;
wire II6560;
wire II6323;
wire II17752;
wire g11599;
wire II5676;
wire II16060;
wire g9920;
wire II5830;
wire II11143;
wire II6924;
wire g10897;
wire II12268;
wire g4511;
wire II14976;
wire II5352;
wire g7431;
wire II6715;
wire g7315;
wire g7285;
wire II15470;
wire g5112;
wire g7497;
wire g7683;
wire g3971;
wire g5813;
wire g10525;
wire g11048;
wire g10930;
wire g8924;
wire g4265;
wire g7732;
wire g2008;
wire II10051;
wire g4920;
wire g5670;
wire g7957;
wire g3055;
wire g5594;
wire g4287;
wire II13554;
wire II6818;
wire II16031;
wire g10769;
wire II14675;
wire g7916;
wire g2563;
wire g6172;
wire g11604;
wire II6572;
wire g11286;
wire g5603;
wire g7140;
wire g4399;
wire II5317;
wire g6621;
wire II16016;
wire g5738;
wire g10356;
wire g2834;
wire g8260;
wire g7344;
wire g11094;
wire g6243;
wire II7600;
wire g9450;
wire g11366;
wire g6468;
wire g7141;
wire g11030;
wire g3473;
wire g11087;
wire g2196;
wire g2067;
wire II7697;
wire g10970;
wire II13773;
wire g2012;
wire g6673;
wire g10646;
wire g8233;
wire II11961;
wire g7362;
wire II14933;
wire g2845;
wire g7145;
wire II14176;
wire g11008;
wire g11346;
wire II16311;
wire g10702;
wire II14405;
wire g9948;
wire g7661;
wire g2751;
wire g8930;
wire g4895;
wire g11543;
wire g7047;
wire g6886;
wire g4941;
wire g7877;
wire g6084;
wire II14534;
wire g10272;
wire II10009;
wire II12568;
wire g10896;
wire II6779;
wire II9362;
wire II5827;
wire g11611;
wire g10386;
wire g10167;
wire II5929;
wire g2272;
wire II16682;
wire II16796;
wire II7034;
wire g6345;
wire II15530;
wire g2229;
wire II15258;
wire g5695;
wire II10514;
wire II9065;
wire g7648;
wire II8877;
wire II11412;
wire g8282;
wire g5260;
wire II5995;
wire g3623;
wire g6329;
wire g5628;
wire g7139;
wire g4501;
wire g7940;
wire g10592;
wire II17525;
wire g10330;
wire g6859;
wire g6287;
wire g10776;
wire g3496;
wire g2405;
wire g7598;
wire g5822;
wire II6962;
wire g11171;
wire II9237;
wire g11403;
wire g7591;
wire g9259;
wire g6863;
wire II17124;
wire II5297;
wire II16286;
wire g9660;
wire g11453;
wire g6521;
wire g7809;
wire II15907;
wire II15691;
wire g9765;
wire g3040;
wire II9165;
wire g4584;
wire g3540;
wire g11262;
wire II13344;
wire g4065;
wire II14272;
wire g4239;
wire II12846;
wire g5757;
wire g5350;
wire g5475;
wire g10827;
wire g8041;
wire II10693;
wire g3769;
wire g10626;
wire g7079;
wire II12939;
wire g4630;
wire g5545;
wire g10746;
wire g5199;
wire g6623;
wire g6184;
wire g5780;
wire g8765;
wire II7330;
wire g8356;
wire g8559;
wire II11262;
wire g4365;
wire II17416;
wire g6681;
wire II11644;
wire g5568;
wire II15347;
wire g4228;
wire g6776;
wire g4491;
wire II14831;
wire g3913;
wire g5279;
wire II15482;
wire g8296;
wire g6179;
wire g7522;
wire g8542;
wire II12126;
wire II9617;
wire g6692;
wire II12153;
wire g9690;
wire II15039;
wire g8444;
wire g9579;
wire g5219;
wire g6056;
wire g5344;
wire g3715;
wire g10900;
wire g6687;
wire g11072;
wire g10907;
wire g10363;
wire g9387;
wire g9669;
wire II13521;
wire g4757;
wire g7769;
wire g8074;
wire g2017;
wire II12186;
wire g10808;
wire g3321;
wire g10079;
wire g4418;
wire II11879;
wire g2132;
wire g11333;
wire g9342;
wire II10966;
wire II5013;
wire g4354;
wire g9652;
wire II6469;
wire g9269;
wire g7930;
wire g7101;
wire II14397;
wire g10558;
wire II9040;
wire II15476;
wire g5521;
wire g7038;
wire g10597;
wire II6330;
wire g11518;
wire II10920;
wire g4379;
wire II12380;
wire g3622;
wire II16264;
wire II17400;
wire II16088;
wire g4617;
wire g5734;
wire II13013;
wire II10030;
wire g7939;
wire g6533;
wire g6190;
wire g4123;
wire g11100;
wire g10136;
wire g4724;
wire II14822;
wire g9934;
wire g2525;
wire g3407;
wire g2242;
wire g5993;
wire II15072;
wire g5824;
wire g8225;
wire g5262;
wire g3334;
wire g4187;
wire g6657;
wire II7002;
wire II8889;
wire g5422;
wire II13403;
wire g7351;
wire g11594;
wire g8102;
wire II7923;
wire g9741;
wire g5744;
wire g11513;
wire g6645;
wire g3628;
wire g6984;
wire g5576;
wire II5913;
wire g8448;
wire g8364;
wire g2060;
wire g6023;
wire II6019;
wire II12592;
wire g4001;
wire g9264;
wire g8722;
wire g6400;
wire g4305;
wire g9821;
wire g9883;
wire II11995;
wire g7430;
wire g6316;
wire g9608;
wire g7211;
wire g6635;
wire II10888;
wire II10520;
wire g6957;
wire g10562;
wire II17240;
wire g7044;
wire g6555;
wire g2753;
wire II13233;
wire II7414;
wire g10104;
wire g4838;
wire g7671;
wire II15900;
wire g7949;
wire II13301;
wire g7097;
wire g6280;
wire g5698;
wire g4420;
wire g3533;
wire g10173;
wire g6877;
wire II17419;
wire g6480;
wire II10024;
wire g10039;
wire g2852;
wire g8742;
wire II10117;
wire II4972;
wire g7601;
wire II6772;
wire g11351;
wire g9714;
wire g9331;
wire g4543;
wire II11306;
wire g10375;
wire II13421;
wire II14645;
wire g2824;
wire g3287;
wire g7065;
wire II13131;
wire II13478;
wire g3433;
wire II14776;
wire II15467;
wire II9159;
wire g10192;
wire g4393;
wire g9726;
wire g8325;
wire g7983;
wire II9007;
wire g10369;
wire II13351;
wire II11602;
wire II15510;
wire g5417;
wire II17231;
wire g9508;
wire g4760;
wire g7625;
wire II7906;
wire II6938;
wire II12145;
wire II6806;
wire g6567;
wire g8097;
wire g10887;
wire II12242;
wire g7779;
wire g10480;
wire II11929;
wire g3365;
wire II8265;
wire II15890;
wire II7931;
wire g2578;
wire II6176;
wire II11201;
wire g7988;
wire g6076;
wire g11559;
wire g4959;
wire II10108;
wire g11213;
wire II13294;
wire g4341;
wire g9945;
wire g8549;
wire II5909;
wire g9867;
wire g11246;
wire g5497;
wire g3274;
wire II5604;
wire g9888;
wire g8303;
wire II7630;
wire II5363;
wire g7221;
wire g7802;
wire g2812;
wire g5768;
wire g6562;
wire g7743;
wire II13397;
wire g5684;
wire g5067;
wire g3267;
wire g2220;
wire II10770;
wire II12779;
wire g8430;
wire g7313;
wire II14133;
wire g4310;
wire g6550;
wire II11882;
wire II13583;
wire g8158;
wire g5856;
wire g8067;
wire g8241;
wire g8575;
wire II5725;
wire II14210;
wire g8478;
wire g6215;
wire g10296;
wire II12694;
wire II13076;
wire g6499;
wire g7567;
wire II10671;
wire g2090;
wire II11629;
wire g11202;
wire g11391;
wire II8815;
wire g3682;
wire g8443;
wire g5223;
wire g4334;
wire g3422;
wire g6619;
wire g3272;
wire g9107;
wire g8595;
wire II16086;
wire g8875;
wire g2516;
wire g6914;
wire II14421;
wire II5565;
wire g8798;
wire II17516;
wire II12093;
wire II13091;
wire II10566;
wire g2569;
wire g8348;
wire g3523;
wire g11338;
wire II15157;
wire II15616;
wire g7119;
wire II17672;
wire g10262;
wire g7547;
wire g11436;
wire g5704;
wire II5251;
wire g10468;
wire g7632;
wire II17494;
wire g3970;
wire g11182;
wire g6910;
wire g8778;
wire g3771;
wire g2117;
wire g6809;
wire g4058;
wire g6716;
wire g3391;
wire g2420;
wire II6403;
wire II8811;
wire II16101;
wire g8820;
wire g8784;
wire g8529;
wire g4550;
wire II17486;
wire g10785;
wire g7402;
wire g7425;
wire g4537;
wire g11442;
wire II11953;
wire g10725;
wire g11272;
wire g2803;
wire g5849;
wire g7082;
wire g5653;
wire g8803;
wire g4453;
wire g5287;
wire II14967;
wire g22;
wire II7612;
wire g8275;
wire g10583;
wire g11487;
wire II9446;
wire II17155;
wire II15639;
wire II15609;
wire II5424;
wire g4515;
wire g2790;
wire II4876;
wire II6881;
wire g6126;
wire g8249;
wire II9734;
wire g4802;
wire g4258;
wire g11254;
wire g3662;
wire g9774;
wire II9826;
wire g6451;
wire g8712;
wire g11057;
wire II15199;
wire g11287;
wire g7054;
wire g10145;
wire g8758;
wire II8786;
wire g2267;
wire g8477;
wire II15795;
wire II9216;
wire g4970;
wire g3093;
wire II7864;
wire g8046;
wire g4489;
wire g5618;
wire g2539;
wire g7826;
wire g3505;
wire g11464;
wire g4639;
wire g4326;
wire g5390;
wire g8671;
wire g10183;
wire II14326;
wire g2713;
wire II15079;
wire g9429;
wire g2085;
wire g2962;
wire g8613;
wire II7840;
wire g10473;
wire II15507;
wire g10394;
wire g3138;
wire g7395;
wire II5858;
wire II14355;
wire g9842;
wire g6708;
wire g5200;
wire II8089;
wire II9564;
wire II12214;
wire II16546;
wire g10715;
wire II16574;
wire II5530;
wire II6199;
wire II12138;
wire II12445;
wire II12867;
wire g5084;
wire II17289;
wire II16589;
wire II10325;
wire II9329;
wire g4480;
wire II6654;
wire g9676;
wire g3328;
wire g6513;
wire g7750;
wire II12171;
wire II12451;
wire II10531;
wire g4572;
wire g2345;
wire g7999;
wire g8343;
wire g9893;
wire g4784;
wire g10253;
wire II9695;
wire g7904;
wire II11280;
wire II6428;
wire g9871;
wire g11644;
wire II16187;
wire II13514;
wire g5232;
wire II11889;
wire II5044;
wire g10498;
wire g6938;
wire II9731;
wire g5192;
wire II11333;
wire g6789;
wire II8551;
wire II5047;
wire II12289;
wire g8176;
wire g8738;
wire II7348;
wire g11657;
wire g5641;
wire g10481;
wire g10469;
wire II11222;
wire II9229;
wire II16580;
wire g5840;
wire g7724;
wire g10451;
wire II13978;
wire g10619;
wire g4567;
wire g9670;
wire g11629;
wire II11821;
wire II16307;
wire g7816;
wire g10752;
wire g7329;
wire g6241;
wire g8755;
wire g5127;
wire g2437;
wire g11186;
wire g1980;
wire g2742;
wire g5837;
wire g2165;
wire g6752;
wire g8570;
wire g2988;
wire II13326;
wire g4881;
wire g10522;
wire II7216;
wire II6043;
wire II11242;
wire g8605;
wire II9574;
wire II5067;
wire g11406;
wire II8259;
wire g10239;
wire g11446;
wire g5528;
wire g5078;
wire g11425;
wire g8185;
wire II5165;
wire g3982;
wire II12397;
wire II7009;
wire II9842;
wire g2099;
wire g2994;
wire g8719;
wire g5397;
wire II8147;
wire g3816;
wire g11015;
wire II11459;
wire II6097;
wire II10286;
wire g6797;
wire g7051;
wire g2391;
wire g10206;
wire g8161;
wire II7886;
wire g4466;
wire g4295;
wire g5172;
wire II6702;
wire g2562;
wire II5089;
wire g7785;
wire g6238;
wire g8629;
wire g3260;
wire g6790;
wire g4204;
wire II11509;
wire g3359;
wire g3104;
wire g7685;
wire g2797;
wire g97;
wire g5912;
wire g7783;
wire g4737;
wire g7389;
wire II11967;
wire II10352;
wire II14127;
wire II13265;
wire g4816;
wire g6713;
wire g5360;
wire g2206;
wire g7686;
wire g6807;
wire g7955;
wire II16781;
wire g2198;
wire g10712;
wire II15811;
wire g5672;
wire II16739;
wire g9348;
wire II7858;
wire g11409;
wire g9647;
wire g10533;
wire g8350;
wire g5605;
wire g8289;
wire II7096;
wire g8659;
wire II9863;
wire g6646;
wire g10110;
wire II6807;
wire II12604;
wire g2479;
wire g11143;
wire II11477;
wire II9581;
wire g2860;
wire g7470;
wire g11075;
wire II10367;
wire g7596;
wire II11122;
wire g5520;
wire g6888;
wire g3708;
wire II12541;
wire II17528;
wire II11695;
wire II16496;
wire II13834;
wire g11480;
wire g10380;
wire g7663;
wire g2531;
wire g3995;
wire g10591;
wire g2215;
wire II14668;
wire g5248;
wire g10700;
wire g2256;
wire g9534;
wire g7751;
wire g6695;
wire g7560;
wire g2219;
wire II9287;
wire II14105;
wire g7772;
wire g4289;
wire II16066;
wire g10251;
wire II5073;
wire g6461;
wire g2022;
wire II16790;
wire g2987;
wire II12384;
wire II17546;
wire II14858;
wire g5033;
wire II12190;
wire g2338;
wire g8421;
wire g3999;
wire II14242;
wire g4316;
wire II11232;
wire g11041;
wire II14367;
wire II11704;
wire g3419;
wire II14257;
wire II9117;
wire g7918;
wire II12300;
wire g2061;
wire II5343;
wire II16024;
wire II17277;
wire II16121;
wire g3097;
wire g8612;
wire II5561;
wire g11197;
wire g5500;
wire II10521;
wire g2538;
wire g7543;
wire II17255;
wire g7890;
wire g8290;
wire g6707;
wire g5890;
wire g2161;
wire g11176;
wire II4883;
wire II13876;
wire g11291;
wire II13454;
wire g2556;
wire g6469;
wire g5708;
wire II4987;
wire g10642;
wire II14010;
wire g8214;
wire II15898;
wire g6639;
wire g7465;
wire g3737;
wire g2331;
wire g8655;
wire II12762;
wire g7823;
wire g6775;
wire g5224;
wire g6170;
wire II16586;
wire g6116;
wire II8663;
wire II7284;
wire g10101;
wire g8390;
wire g8377;
wire g11086;
wire g10890;
wire II12318;
wire II4973;
wire g8774;
wire g9747;
wire g5723;
wire II6714;
wire g11347;
wire g5031;
wire g7792;
wire g8737;
wire g10850;
wire g4263;
wire g5509;
wire g4336;
wire g8966;
wire II10759;
wire II15296;
wire g6324;
wire g4426;
wire g3625;
wire g2131;
wire g4912;
wire II11085;
wire g9415;
wire II14239;
wire g9720;
wire II5626;
wire II17213;
wire g7540;
wire II5284;
wire g9845;
wire g7259;
wire g4081;
wire II11942;
wire g3907;
wire g10425;
wire II7946;
wire g6127;
wire II7396;
wire II16604;
wire g10549;
wire II6074;
wire g4538;
wire g4788;
wire g5094;
wire g5263;
wire II10952;
wire g7184;
wire II6504;
wire II6233;
wire g3460;
wire g5241;
wire g4514;
wire II10932;
wire g11278;
wire II12589;
wire g5825;
wire g9192;
wire II11420;
wire II8506;
wire II11653;
wire II8123;
wire g10190;
wire II17302;
wire II11936;
wire II6947;
wire g11148;
wire g3813;
wire g4592;
wire g3812;
wire g7303;
wire g11539;
wire II15338;
wire g9025;
wire g11320;
wire g11416;
wire II14204;
wire g10056;
wire g4250;
wire II11049;
wire g8626;
wire g2644;
wire g6802;
wire II16214;
wire g4521;
wire g9698;
wire g8173;
wire II12499;
wire II10706;
wire II7729;
wire g9782;
wire g8336;
wire g6038;
wire II8640;
wire g6288;
wire II6789;
wire g1965;
wire g3545;
wire g9519;
wire II12056;
wire II7659;
wire II13445;
wire g11637;
wire g10799;
wire II15694;
wire II14678;
wire II5070;
wire II7118;
wire II13258;
wire g10051;
wire g4217;
wire g3753;
wire g6624;
wire g11265;
wire g9703;
wire g5886;
wire g6315;
wire II13952;
wire II10861;
wire g5639;
wire II8324;
wire g3940;
wire g8236;
wire II12223;
wire g5482;
wire II9776;
wire g7438;
wire II16676;
wire g5569;
wire g5107;
wire g7334;
wire g3942;
wire II13489;
wire g3967;
wire II14119;
wire II5516;
wire g6019;
wire g8359;
wire g10169;
wire II9857;
wire g2825;
wire g11605;
wire g8416;
wire g3520;
wire g11209;
wire g6443;
wire g4766;
wire II4966;
wire g9725;
wire g11646;
wire II14217;
wire II5410;
wire g3978;
wire g8451;
wire g6582;
wire g6432;
wire g4739;
wire g11309;
wire II9433;
wire g4878;
wire g6904;
wire g9813;
wire g5917;
wire g10244;
wire g4113;
wire g11229;
wire g8147;
wire II5311;
wire II12159;
wire g10579;
wire g4339;
wire g6964;
wire II13354;
wire g6560;
wire II17265;
wire g8439;
wire g5116;
wire g9642;
wire g2623;
wire II12793;
wire II8911;
wire g10886;
wire II14531;
wire g10658;
wire II15870;
wire g10932;
wire g8195;
wire II13990;
wire g10121;
wire II14970;
wire g2176;
wire II7636;
wire g9658;
wire g4141;
wire II11632;
wire II6805;
wire g2507;
wire g11475;
wire g2890;
wire g9966;
wire II8024;
wire g9864;
wire II6510;
wire II4954;
wire II14485;
wire g8089;
wire II12627;
wire g7929;
wire g4050;
wire g10317;
wire g5416;
wire II9575;
wire II5605;
wire g3790;
wire g6875;
wire II13285;
wire g8514;
wire g9803;
wire g8265;
wire g7574;
wire II16799;
wire g11463;
wire g2854;
wire g11288;
wire g11152;
wire II17318;
wire g11212;
wire g6341;
wire g11096;
wire g10432;
wire II15193;
wire g5299;
wire II13017;
wire g10676;
wire II17552;
wire II10927;
wire g10876;
wire II16638;
wire g4893;
wire II12282;
wire g5677;
wire II12838;
wire II8253;
wire g6274;
wire g8284;
wire g7232;
wire g6247;
wire II11566;
wire g6728;
wire II5893;
wire g9817;
wire g5100;
wire II6220;
wire g1975;
wire g5182;
wire g7692;
wire II15209;
wire g5731;
wire II10607;
wire g6816;
wire g8127;
wire g10087;
wire II11686;
wire g11097;
wire II11094;
wire g8812;
wire g7651;
wire II13245;
wire II8848;
wire II6356;
wire II9141;
wire g4934;
wire II6580;
wire g5613;
wire g2344;
wire II7820;
wire II4929;
wire g8649;
wire II11800;
wire II8717;
wire g2270;
wire II11975;
wire g8729;
wire g4490;
wire g5841;
wire II8228;
wire g2677;
wire g3037;
wire g10974;
wire g5029;
wire g9838;
wire g4499;
wire g3246;
wire g2940;
wire II16196;
wire II10201;
wire g7619;
wire g3860;
wire II6080;
wire II11348;
wire g3112;
wire g10735;
wire II13320;
wire g9613;
wire g6832;
wire g11654;
wire g4272;
wire II5438;
wire II12400;
wire II12032;
wire g6031;
wire g5772;
wire g10138;
wire II11537;
wire II14709;
wire g7519;
wire g10439;
wire II13645;
wire II16200;
wire g5189;
wire II15190;
wire II17733;
wire g8730;
wire g3938;
wire g5818;
wire II15526;
wire II12062;
wire g5286;
wire g4671;
wire g2056;
wire g7780;
wire II17500;
wire II11790;
wire g4820;
wire II14444;
wire II6976;
wire g8878;
wire II12412;
wire II6676;
wire II9525;
wire g10401;
wire g2500;
wire g11433;
wire g4827;
wire g8868;
wire g11220;
wire g10540;
wire II13918;
wire g8109;
wire II12430;
wire g6296;
wire g7846;
wire II12409;
wire g7009;
wire II9620;
wire II4948;
wire g11028;
wire II5658;
wire g3878;
wire g2757;
wire g5719;
wire II9171;
wire II13618;
wire g6846;
wire II9965;
wire g8329;
wire g3758;
wire g8505;
wire II6111;
wire g2945;
wire g6137;
wire g8708;
wire g2046;
wire g9828;
wire II17158;
wire g6347;
wire II13370;
wire II16458;
wire g10080;
wire g6003;
wire II11590;
wire g10564;
wire II11677;
wire g10234;
wire g6485;
wire g6412;
wire g6385;
wire g9593;
wire g3705;
wire II9105;
wire II8625;
wire g11496;
wire g8934;
wire II13504;
wire g6332;
wire g5314;
wire II5388;
wire II8237;
wire II15617;
wire g9911;
wire g3207;
wire II8462;
wire g8003;
wire g7573;
wire g8140;
wire g10478;
wire g8157;
wire II5366;
wire II15320;
wire g7581;
wire g7532;
wire g4713;
wire II6661;
wire g7443;
wire g9413;
wire g2911;
wire g9661;
wire g5145;
wire g5811;
wire II10018;
wire II6520;
wire g11413;
wire g7510;
wire II7763;
wire g7189;
wire g10865;
wire g8560;
wire g11150;
wire g6145;
wire g7584;
wire g10745;
wire g7966;
wire g4465;
wire g7394;
wire g5664;
wire g6122;
wire g8014;
wire g7959;
wire g3723;
wire II7300;
wire g4164;
wire II12577;
wire g8254;
wire II9557;
wire g8881;
wire II9947;
wire g10696;
wire g9995;
wire II13806;
wire g5779;
wire g11107;
wire g8274;
wire g8267;
wire g3799;
wire g5934;
wire II11011;
wire II7438;
wire g9734;
wire g10325;
wire g6546;
wire g10670;
wire g8297;
wire g7631;
wire g6733;
wire g3389;
wire g6758;
wire g3011;
wire g6531;
wire g7767;
wire g2316;
wire g9586;
wire g3719;
wire II5468;
wire II10739;
wire g8388;
wire II16817;
wire g2006;
wire II8575;
wire g8839;
wire g7853;
wire g8697;
wire g8150;
wire g7886;
wire g7256;
wire II4912;
wire g8552;
wire II9851;
wire g7502;
wire g10452;
wire II16073;
wire g8714;
wire II10630;
wire g6306;
wire g7293;
wire g10433;
wire g2872;
wire II9839;
wire g11435;
wire g6709;
wire II9213;
wire II7509;
wire g2506;
wire g2350;
wire g6580;
wire II8315;
wire g10818;
wire g4013;
wire g2227;
wire g2209;
wire II14443;
wire g10063;
wire g11404;
wire g7741;
wire II9845;
wire II6914;
wire g7722;
wire II11450;
wire g10392;
wire II10843;
wire g5174;
wire g11452;
wire g11443;
wire g4905;
wire II11935;
wire g4906;
wire II12136;
wire g6826;
wire g5859;
wire II9377;
wire g8573;
wire g6318;
wire g4993;
wire g7697;
wire g4463;
wire g10075;
wire II11970;
wire g6337;
wire II7668;
wire II5221;
wire g3776;
wire g9856;
wire g10860;
wire II15048;
wire g11203;
wire g4298;
wire g8635;
wire II14561;
wire g4541;
wire g8828;
wire II10620;
wire II9224;
wire II17410;
wire g3041;
wire g8234;
wire g6912;
wire II6287;
wire g7374;
wire g5121;
wire g6515;
wire II6447;
wire g9427;
wire g7710;
wire g7050;
wire g11579;
wire g2763;
wire g10032;
wire g5839;
wire g11183;
wire II14546;
wire g7076;
wire II14249;
wire g10682;
wire g3373;
wire g6425;
wire g4003;
wire g8180;
wire g8379;
wire g5643;
wire g11244;
wire II9519;
wire II7766;
wire g6854;
wire g4762;
wire g8694;
wire g8272;
wire g10305;
wire g10227;
wire II16298;
wire g11380;
wire g11627;
wire II5579;
wire g11582;
wire II17170;
wire II9923;
wire II9602;
wire g6724;
wire g7287;
wire g8252;
wire g5592;
wire g7909;
wire g3717;
wire g10867;
wire g3988;
wire II11021;
wire g4785;
wire II6747;
wire II6837;
wire II8234;
wire II6778;
wire g6927;
wire II17179;
wire g2322;
wire g10359;
wire g5751;
wire g7125;
wire g6787;
wire g3392;
wire g5903;
wire g10718;
wire g7033;
wire II7333;
wire II6624;
wire II9860;
wire g10574;
wire g7368;
wire II11249;
wire II6091;
wire II11278;
wire II10012;
wire g4746;
wire II8080;
wire g9555;
wire g2903;
wire g9088;
wire gbuf11;
wire II10756;
wire g4486;
wire g2814;
wire g5735;
wire g10635;
wire II5837;
wire g6407;
wire II6144;
wire g8060;
wire g7361;
wire II17356;
wire g8043;
wire g11415;
wire g6166;
wire g7265;
wire II5805;
wire g5510;
wire II9394;
wire g3424;
wire g2034;
wire II8011;
wire g4203;
wire II8490;
wire g2517;
wire g5118;
wire II17435;
wire g6906;
wire II12638;
wire g4270;
wire g4185;
wire II14077;
wire g2877;
wire g2510;
wire g8873;
wire g8184;
wire II17441;
wire g2238;
wire g11372;
wire g6834;
wire II11540;
wire g2799;
wire g7961;
wire g10290;
wire II11810;
wire II10503;
wire g11279;
wire II10682;
wire g7353;
wire II7351;
wire g1994;
wire II8139;
wire g2804;
wire g8794;
wire g5205;
wire g4582;
wire II5677;
wire II14499;
wire g9617;
wire g6105;
wire g4577;
wire g5398;
wire g11281;
wire II13039;
wire II6880;
wire g6058;
wire g9897;
wire II12610;
wire g8786;
wire g2234;
wire II5127;
wire g4476;
wire g9957;
wire II15308;
wire g7920;
wire g11598;
wire g11459;
wire g11393;
wire g2121;
wire II13439;
wire g9312;
wire g7346;
wire g10261;
wire g2269;
wire g6448;
wire II15269;
wire II8499;
wire g2896;
wire g10424;
wire II9323;
wire II10258;
wire g10207;
wire g11055;
wire g7459;
wire II11898;
wire g5523;
wire II5649;
wire g5620;
wire g8322;
wire g8345;
wire II16667;
wire g3271;
wire g8745;
wire g10554;
wire g5851;
wire g5742;
wire g10899;
wire g5502;
wire g7036;
wire II5263;
wire II8278;
wire g5027;
wire II17739;
wire g2557;
wire g4590;
wire II5599;
wire g5705;
wire g5808;
wire II16169;
wire g5091;
wire g8810;
wire g7927;
wire II11100;
wire g5651;
wire g6573;
wire g3664;
wire g3500;
wire g9891;
wire II17206;
wire II9956;
wire II7456;
wire g11065;
wire II16484;
wire II9505;
wire g5800;
wire g8476;
wire g9922;
wire II11269;
wire II12286;
wire g2792;
wire g4533;
wire g9929;
wire g9390;
wire g7719;
wire g6919;
wire II5041;
wire g6430;
wire g11397;
wire II6143;
wire II16500;
wire II13128;
wire g4255;
wire II5963;
wire II5427;
wire II6317;
wire g6557;
wire II15583;
wire g9591;
wire g11591;
wire II16610;
wire g7599;
wire g8305;
wire g7607;
wire g2750;
wire g5683;
wire g4950;
wire g6584;
wire g4348;
wire g3543;
wire g6503;
wire II12683;
wire g6041;
wire g11329;
wire II13206;
wire II5164;
wire g11589;
wire g10855;
wire II11725;
wire II8851;
wire g8406;
wire g6793;
wire g4415;
wire g11012;
wire II10984;
wire g4988;
wire g10441;
wire II15749;
wire II7642;
wire g4605;
wire g10289;
wire II17657;
wire g3431;
wire g4831;
wire g4070;
wire II15891;
wire g2005;
wire g10822;
wire II8476;
wire II7151;
wire g8535;
wire II10096;
wire II12783;
wire II9935;
wire II16280;
wire II10846;
wire g6282;
wire g3531;
wire II10828;
wire g2957;
wire g10367;
wire g4589;
wire g9823;
wire g9762;
wire g6641;
wire g7898;
wire II9486;
wire g10162;
wire g10884;
wire g9886;
wire g6051;
wire g8827;
wire g10556;
wire II7176;
wire g5213;
wire II6193;
wire g2336;
wire g8958;
wire g11603;
wire g2107;
wire g7349;
wire g5567;
wire g4184;
wire g10170;
wire g9905;
wire g8843;
wire g6565;
wire g11353;
wire II17713;
wire g4383;
wire g5879;
wire g8723;
wire II5619;
wire II17070;
wire g4718;
wire g10280;
wire g4293;
wire g5267;
wire II11608;
wire II17234;
wire g11019;
wire g10910;
wire II7157;
wire g7776;
wire g8414;
wire g11225;
wire g6264;
wire II6726;
wire II13317;
wire II9090;
wire II16660;
wire II14558;
wire g3363;
wire g5686;
wire g7948;
wire II17584;
wire g7206;
wire g2100;
wire g2979;
wire g8763;
wire II15326;
wire g4522;
wire g7337;
wire g11428;
wire g6861;
wire II12045;
wire g6204;
wire g10372;
wire II9883;
wire g2431;
wire g6971;
wire II6955;
wire II10111;
wire g6894;
wire g5669;
wire g6868;
wire g3164;
wire g5221;
wire g5273;
wire g6939;
wire g4614;
wire II17678;
wire g10768;
wire II7372;
wire g11625;
wire g8606;
wire II10698;
wire II10434;
wire g5999;
wire g8441;
wire g10906;
wire g9654;
wire g9691;
wire II13539;
wire g6177;
wire II10795;
wire g10345;
wire g4370;
wire g9557;
wire g1997;
wire g10362;
wire g6688;
wire g10620;
wire g6131;
wire g7931;
wire g4555;
wire II12559;
wire g10787;
wire g7527;
wire g6097;
wire g4233;
wire gbuf8;
wire II12511;
wire II11109;
wire II6163;
wire II5618;
wire g4192;
wire II10689;
wire II8351;
wire II15229;
wire II13394;
wire g4106;
wire g7986;
wire g2543;
wire II15415;
wire II6388;
wire g11335;
wire g4352;
wire II15632;
wire II12369;
wire g8095;
wire g7308;
wire II12357;
wire g9773;
wire g5473;
wire g6193;
wire g5900;
wire g4391;
wire g6062;
wire g2970;
wire II5612;
wire g9526;
wire g4347;
wire II5296;
wire g3408;
wire II6065;
wire g3762;
wire g2641;
wire g7310;
wire II13959;
wire g4774;
wire II14309;
wire g3071;
wire g5544;
wire g6092;
wire g9853;
wire g3387;
wire II12372;
wire g2564;
wire II5812;
wire g8974;
wire g6590;
wire g8989;
wire g3632;
wire II15172;
wire g4005;
wire g3323;
wire g9576;
wire g5257;
wire II16081;
wire g7217;
wire II11869;
wire g4455;
wire g9861;
wire II15374;
wire II6373;
wire g2088;
wire g5867;
wire g10889;
wire g11293;
wire II15879;
wire II14278;
wire II12180;
wire g5150;
wire g11502;
wire II6068;
wire II12460;
wire g7622;
wire II11778;
wire g8776;
wire g5008;
wire g6069;
wire g11519;
wire II16258;
wire II16145;
wire II16950;
wire g6908;
wire g7301;
wire II15051;
wire g2302;
wire g11466;
wire II17591;
wire g8160;
wire g10596;
wire g9150;
wire g6528;
wire II5840;
wire II16863;
wire g7993;
wire II10412;
wire II8858;
wire g7976;
wire g9881;
wire g9932;
wire II17334;
wire g2451;
wire g8020;
wire II15409;
wire II7420;
wire g6525;
wire g11315;
wire II15536;
wire g9847;
wire g8048;
wire g7814;
wire g5005;
wire g2130;
wire II16537;
wire II5525;
wire g11178;
wire II13560;
wire g8759;
wire g7068;
wire g5082;
wire II7935;
wire g6445;
wire g10276;
wire g11302;
wire II13010;
wire g4437;
wire g6249;
wire g11647;
wire g6756;
wire g8029;
wire g6632;
wire II13530;
wire g4977;
wire g8410;
wire g10446;
wire g11322;
wire II9665;
wire g2642;
wire g6169;
wire g9341;
wire g5626;
wire g2349;
wire g3627;
wire g3462;
wire g8499;
wire g9453;
wire g7638;
wire g3426;
wire II14391;
wire g10797;
wire II13482;
wire II8396;
wire g6700;
wire g5403;
wire II12026;
wire g10655;
wire g6897;
wire g11099;
wire g7182;
wire II6477;
wire g11511;
wire II9191;
wire g5944;
wire g10094;
wire g6237;
wire g4474;
wire II15181;
wire g6080;
wire g7820;
wire g4505;
wire II6343;
wire g4345;
wire II13642;
wire II11515;
wire g11418;
wire g5507;
wire g8209;
wire g8791;
wire g3518;
wire II16632;
wire II9807;
wire II9443;
wire g8700;
wire II11584;
wire II5024;
wire II9308;
wire II12103;
wire II11794;
wire g5480;
wire g2041;
wire II16814;
wire g10312;
wire g5884;
wire II12919;
wire g2649;
wire g8334;
wire g10157;
wire g6800;
wire g6087;
wire g6216;
wire II6187;
wire II10123;
wire g5423;
wire II16001;
wire II11807;
wire II7726;
wire g7332;
wire II7318;
wire g11063;
wire g10267;
wire g2985;
wire g5096;
wire II7800;
wire g8964;
wire II13332;
wire g6036;
wire g5114;
wire g7092;
wire II12813;
wire g10284;
wire g2493;
wire g11552;
wire g9431;
wire g6917;
wire g7380;
wire II8676;
wire g11635;
wire II5034;
wire g3909;
wire g8585;
wire g6674;
wire g2264;
wire g8154;
wire g8971;
wire II5847;
wire II13559;
wire g4424;
wire g7673;
wire II11061;
wire II13283;
wire g7436;
wire g4441;
wire II11916;
wire g8819;
wire g6947;
wire g2120;
wire g4868;
wire II16105;
wire g11640;
wire g7387;
wire g9827;
wire g5899;
wire II12472;
wire g2846;
wire II13624;
wire g7953;
wire g2560;
wire II6812;
wire g2258;
wire g7688;
wire g2395;
wire II10789;
wire g10069;
wire g10040;
wire g2346;
wire II14672;
wire g5535;
wire g2210;
wire g6078;
wire II14494;
wire II16507;
wire g5538;
wire g9205;
wire g7594;
wire g8928;
wire II16366;
wire g3440;
wire g5252;
wire g11421;
wire II5833;
wire II6001;
wire g7902;
wire g10531;
wire II12544;
wire g6648;
wire g7944;
wire II7707;
wire g6303;
wire II13886;
wire II10858;
wire g9645;
wire g10542;
wire g9596;
wire II16938;
wire g2037;
wire g11073;
wire g8419;
wire g10335;
wire g6696;
wire g6575;
wire g9473;
wire g8299;
wire g3060;
wire II7260;
wire g6652;
wire g11174;
wire g11110;
wire g10772;
wire II9273;
wire g6291;
wire g5587;
wire II8514;
wire g1992;
wire II12307;
wire II5460;
wire II9399;
wire g4444;
wire g3087;
wire II14537;
wire g9851;
wire g6760;
wire II14528;
wire II5111;
wire g3997;
wire II17261;
wire g9944;
wire g5168;
wire g11340;
wire g7770;
wire II8180;
wire g2773;
wire g6596;
wire g8568;
wire g5843;
wire g4580;
wire g8006;
wire II15992;
wire g8423;
wire g11349;
wire g2821;
wire g7790;
wire II10370;
wire g5648;
wire II15595;
wire g8752;
wire II15817;
wire g2880;
wire II13117;
wire g6855;
wire g9924;
wire g4269;
wire II4985;
wire II9290;
wire g7130;
wire g2760;
wire g10892;
wire II6395;
wire II10592;
wire g11556;
wire g10343;
wire II12424;
wire g2755;
wire II15704;
wire II8771;
wire g5721;
wire g2862;
wire g7476;
wire g5597;
wire g4389;
wire II14687;
wire g4748;
wire II14473;
wire II15176;
wire g4735;
wire g4078;
wire g4280;
wire g3351;
wire II13666;
wire II6917;
wire g6881;
wire II4978;
wire g10382;
wire g3378;
wire g5615;
wire g2103;
wire g11619;
wire II13030;
wire II4971;
wire g7736;
wire g11083;
wire g4439;
wire g7479;
wire g11652;
wire g3636;
wire II14179;
wire g5590;
wire g2732;
wire g8614;
wire g8178;
wire II11505;
wire g11043;
wire g4290;
wire g10199;
wire g4791;
wire g2251;
wire g5827;
wire g6387;
wire II6690;
wire g7990;
wire II10898;
wire g2076;
wire g7799;
wire g10497;
wire g9601;
wire g5877;
wire g3380;
wire II6907;
wire g7765;
wire II9905;
wire g3306;
wire II7429;
wire II15517;
wire g6452;
wire g8706;
wire g6410;
wire g9967;
wire g5353;
wire g10705;
wire II9652;
wire g8424;
wire g8432;
wire g10538;
wire II16941;
wire g8732;
wire g2163;
wire g2808;
wire g6095;
wire g4996;
wire II14376;
wire g7844;
wire g7703;
wire g11035;
wire II15589;
wire g6661;
wire g6267;
wire g7582;
wire g4099;
wire g8480;
wire g5284;
wire II10189;
wire g4673;
wire II6538;
wire g2502;
wire II11668;
wire II5136;
wire g4142;
wire II11909;
wire II11671;
wire g5790;
wire g5180;
wire II13732;
wire II10946;
wire II12822;
wire II7465;
wire II9150;
wire g4125;
wire II13506;
wire II11650;
wire g10035;
wire g2305;
wire g10131;
wire II5795;
wire g4885;
wire II5713;
wire g5187;
wire II12993;
wire g5784;
wire g9358;
wire g8220;
wire g11159;
wire g7530;
wire II5570;
wire g7964;
wire g10511;
wire g7995;
wire g5730;
wire g8386;
wire II13678;
wire II9188;
wire g4367;
wire g9588;
wire g8120;
wire g11618;
wire g2217;
wire g6353;
wire g6735;
wire g7981;
wire g6983;
wire II4910;
wire II16479;
wire II16595;
wire II15427;
wire II11166;
wire g7524;
wire II8973;
wire g2947;
wire II8642;
wire g11504;
wire II7017;
wire g8155;
wire g7504;
wire g5862;
wire g4241;
wire II8577;
wire g2201;
wire g9694;
wire g7187;
wire g10323;
wire g6120;
wire gbuf1;
wire II4786;
wire g8269;
wire g8547;
wire II6671;
wire g11235;
wire g9258;
wire g10672;
wire g7851;
wire g4313;
wire g7445;
wire II5998;
wire g4963;
wire II15744;
wire g2055;
wire g2952;
wire g5795;
wire g10690;
wire g7034;
wire g9010;
wire II15717;
wire II12150;
wire II9598;
wire g3766;
wire g11439;
wire g5701;
wire g8135;
wire g5484;
wire g11399;
wire g3937;
wire g8169;
wire II6367;
wire g11337;
wire g10236;
wire g4711;
wire g1991;
wire g2436;
wire II13255;
wire g8739;
wire g5270;
wire g8888;
wire g3103;
wire g7273;
wire g9917;
wire II6738;
wire II4820;
wire g4105;
wire II14055;
wire g9993;
wire g3226;
wire g10256;
wire II13941;
wire g7225;
wire g4449;
wire g11227;
wire g4775;
wire g3110;
wire g5770;
wire II10541;
wire II12496;
wire g2240;
wire II4964;
wire g5300;
wire II16217;
wire g7545;
wire g6149;
wire II12174;
wire II12053;
wire II5325;
wire g8311;
wire g7134;
wire g7291;
wire II6077;
wire II7677;
wire g9723;
wire II17305;
wire II8164;
wire g10228;
wire II7564;
wire g11577;
wire II13837;
wire g7558;
wire II10293;
wire g10766;
wire g7758;
wire II6733;
wire g8463;
wire II5224;
wire II17104;
wire g6273;
wire g6814;
wire g2639;
wire II7223;
wire II17249;
wire g5739;
wire g8948;
wire II13992;
wire II16038;
wire II10885;
wire g11026;
wire II11543;
wire II14452;
wire g7557;
wire II14123;
wire g5919;
wire g2748;
wire II11152;
wire g4296;
wire g10243;
wire g10492;
wire g4231;
wire g6339;
wire g8571;
wire g5941;
wire II14083;
wire g10315;
wire g11561;
wire II7875;
wire g3222;
wire g8464;
wire g10674;
wire g6278;
wire g5666;
wire II10589;
wire II16289;
wire II15219;
wire II13236;
wire g6103;
wire g4781;
wire II16461;
wire II5002;
wire II11973;
wire g9532;
wire g6343;
wire g4331;
wire g7660;
wire II9946;
wire II6443;
wire g4214;
wire g2963;
wire g2828;
wire g8263;
wire g4167;
wire gbuf6;
wire g10936;
wire g3976;
wire g6054;
wire g9615;
wire g4279;
wire II15441;
wire g6001;
wire g10200;
wire g10248;
wire g3695;
wire g10852;
wire g8145;
wire II13242;
wire g2778;
wire g8939;
wire g6874;
wire g2194;
wire g4458;
wire g6254;
wire g11587;
wire II16468;
wire II4920;
wire g4726;
wire II4935;
wire II5878;
wire II9135;
wire g10484;
wire g9490;
wire g8125;
wire g10128;
wire g7103;
wire g10874;
wire g7617;
wire g2801;
wire g10665;
wire g6540;
wire g6570;
wire g9941;
wire g3370;
wire g10733;
wire II9415;
wire g10759;
wire g8104;
wire g7413;
wire g4083;
wire g9292;
wire g2173;
wire II10553;
wire II10891;
wire g11473;
wire g4876;
wire g6071;
wire II5478;
wire II15787;
wire II12601;
wire g3863;
wire g8409;
wire g3039;
wire g9815;
wire g4497;
wire g5089;
wire g5109;
wire g2353;
wire II11617;
wire g7375;
wire g5104;
wire g11447;
wire g11205;
wire g4807;
wire g7748;
wire g5425;
wire g7406;
wire g3485;
wire g4323;
wire II15983;
wire II11572;
wire g5633;
wire g9103;
wire II9833;
wire g8473;
wire II8678;
wire II7710;
wire g10292;
wire II8268;
wire g2965;
wire g2873;
wire g8871;
wire g10934;
wire II6138;
wire II13188;
wire g4318;
wire g6836;
wire II7513;
wire g4007;
wire g6667;
wire II12878;
wire g7325;
wire II11146;
wire g7004;
wire g10299;
wire II7210;
wire g7924;
wire g11253;
wire II13909;
wire II7363;
wire g4376;
wire g8251;
wire g5853;
wire II9123;
wire g2070;
wire g6164;
wire II10156;
wire II7732;
wire g2081;
wire g11023;
wire g8435;
wire g10862;
wire II6424;
wire g4767;
wire g3318;
wire g10513;
wire g6552;
wire g10820;
wire g11223;
wire g9079;
wire II17447;
wire g7922;
wire g1962;
wire II12930;
wire II7757;
wire II10804;
wire II13307;
wire g5573;
wire g11623;
wire II14519;
wire g8816;
wire g5619;
wire g10202;
wire II7462;
wire g6245;
wire g4562;
wire II17438;
wire II6799;
wire g8743;
wire g8320;
wire g10422;
wire g9778;
wire g6702;
wire II12265;
wire II14130;
wire II12439;
wire g3205;
wire g6934;
wire g4253;
wire II8885;
wire II11981;
wire g2299;
wire II6771;
wire g10429;
wire II7387;
wire g3413;
wire g10728;
wire g4201;
wire g11395;
wire g7258;
wire g4535;
wire g8825;
wire II10192;
wire g5802;
wire g7421;
wire g2960;
wire II5886;
wire g9959;
wire II17384;
wire II12532;
wire g9522;
wire g4088;
wire g9528;
wire g8955;
wire II9612;
wire g4518;
wire g9411;
wire g7717;
wire II11623;
wire g7612;
wire g8474;
wire g2655;
wire g10487;
wire II14585;
wire g9899;
wire II5265;
wire II16178;
wire g8182;
wire g2794;
wire g6256;
wire g2236;
wire g4209;
wire g5688;
wire g9854;
wire g3331;
wire g7127;
wire g10390;
wire II13561;
wire g10143;
wire II8116;
wire g7123;
wire g10707;
wire g4721;
wire g11165;
wire g5645;
wire II15278;
wire II6616;
wire g9671;
wire g7720;
wire II11211;
wire II8989;
wire g5043;
wire g3730;
wire g11608;
wire g8482;
wire II10437;
wire g11258;
wire g6718;
wire g2225;
wire II14793;
wire g4052;
wire g4073;
wire II11338;
wire g2180;
wire II14109;
wire g6537;
wire g4011;
wire g7788;
wire II5593;
wire g7738;
wire g11548;
wire II16644;
wire g5123;
wire g8079;
wire II11956;
wire II9699;
wire g5789;
wire g6517;
wire g10608;
wire g2765;
wire g9553;
wire g6325;
wire II7236;
wire g6046;
wire g10271;
wire g8771;
wire g8617;
wire II11005;
wire II13803;
wire g8008;
wire g5419;
wire g6423;
wire g9353;
wire g5902;
wire g10680;
wire g11318;
wire II15448;
wire II5854;
wire g7705;
wire II14805;
wire II14385;
wire II12274;
wire II14955;
wire II6921;
wire g4368;
wire g6113;
wire II10535;
wire II12165;
wire II7339;
wire II14209;
wire g5126;
wire II11447;
wire g2094;
wire II16255;
wire II13900;
wire g7880;
wire g4891;
wire g11622;
wire g8601;
wire gbuf13;
wire g2186;
wire g4325;
wire II12514;
wire II9311;
wire g5691;
wire g5896;
wire II13068;
wire g7340;
wire g5674;
wire II8545;
wire II10477;
wire g7366;
wire II12113;
wire g7220;
wire g5679;
wire II8487;
wire g6711;
wire g10552;
wire g7059;
wire g6470;
wire g5236;
wire g4484;
wire g7322;
wire g2232;
wire II10710;
wire g3263;
wire g7204;
wire g2998;
wire g7271;
wire g1984;
wire g5176;
wire g7727;
wire II16052;
wire II5620;
wire g11481;
wire g7319;
wire g4261;
wire g8608;
wire g7031;
wire g10435;
wire II15559;
wire II9571;
wire g4243;
wire g4618;
wire II12261;
wire II15431;
wire g4198;
wire II5818;
wire g2433;
wire g10716;
wire II7776;
wire II6988;
wire II8211;
wire II15520;
wire II17684;
wire g11478;
wire g11157;
wire g10303;
wire g11468;
wire II15383;
wire g8625;
wire g4903;
wire II10971;
wire II9813;
wire g5997;
wire g3764;
wire g9711;
wire II12454;
wire II13659;
wire g10803;
wire g9656;
wire g7900;
wire g7040;
wire g5073;
wire II11351;
wire g7805;
wire g9663;
wire g10443;
wire g10904;
wire g2837;
wire II9111;
wire g8769;
wire g6026;
wire g5753;
wire g8100;
wire II17353;
wire g2789;
wire II15287;
wire II9205;
wire g9563;
wire II11322;
wire II6990;
wire g3015;
wire II11360;
wire g3255;
wire II13537;
wire g7946;
wire II14116;
wire g6547;
wire g6235;
wire II12232;
wire g3819;
wire g9771;
wire g9757;
wire g4728;
wire g2480;
wire II8290;
wire g9761;
wire II10066;
wire g6060;
wire g6990;
wire g7463;
wire g9990;
wire II10456;
wire II13888;
wire g8200;
wire g9731;
wire g10360;
wire g4121;
wire g10622;
wire g10600;
wire g7933;
wire g5469;
wire g8961;
wire II5866;
wire g4969;
wire g6502;
wire g8190;
wire II17271;
wire g8733;
wire g7629;
wire g5275;
wire g8099;
wire g4495;
wire II10907;
wire g5542;
wire g4359;
wire g5720;
wire g8546;
wire g4235;
wire g6194;
wire g11457;
wire g8553;
wire g11242;
wire g7355;
wire g2910;
wire II15473;
wire g9256;
wire g9960;
wire II11824;
wire II11528;
wire g10187;
wire II15485;
wire g3536;
wire g11146;
wire II7956;
wire II11464;
wire g5254;
wire g8886;
wire g2110;
wire II12953;
wire g7590;
wire g10411;
wire g5471;
wire g8218;
wire II8900;
wire g8050;
wire II8250;
wire g9265;
wire g8987;
wire g2529;
wire g6950;
wire g5401;
wire g6067;
wire II12092;
wire g7978;
wire g3634;
wire II16650;
wire g10352;
wire II6126;
wire II5372;
wire II5210;
wire g11307;
wire g10901;
wire II14555;
wire II12293;
wire g3428;
wire g7624;
wire g10389;
wire g11053;
wire g10780;
wire II12074;
wire g6626;
wire g7812;
wire II8527;
wire g5555;
wire g9938;
wire g11498;
wire II14910;
wire II9388;
wire II6016;
wire g2245;
wire II5584;
wire II13592;
wire g9930;
wire g9768;
wire g10047;
wire g9507;
wire g6943;
wire II8520;
wire II6630;
wire g7025;
wire II4780;
wire g6586;
wire II5142;
wire g9425;
wire g7106;
wire II16626;
wire II12099;
wire g8039;
wire g4753;
wire g8229;
wire g11218;
wire II6224;
wire g6090;
wire II15864;
wire II9792;
wire II17371;
wire II10093;
wire II5765;
wire g7605;
wire II11252;
wire g7822;
wire g4952;
wire g7416;
wire II16772;
wire g3621;
wire g4361;
wire II10648;
wire g2885;
wire g7209;
wire g8193;
wire g7350;
wire g10387;
wire II13191;
wire g10185;
wire g11426;
wire g2381;
wire II15965;
wire II10033;
wire g6220;
wire g4300;
wire II6557;
wire g5718;
wire II10904;
wire II15698;
wire II9320;
wire II10724;
wire g8115;
wire g8360;
wire g4770;
wire II8036;
wire g7074;
wire g10774;
wire g5420;
wire g3345;
wire g10687;
wire g5349;
wire II11345;
wire g6479;
wire g11450;
wire g6509;
wire II5966;
wire g2101;
wire g5727;
wire II6932;
wire II17755;
wire g5470;
wire g7516;
wire g10577;
wire II8429;
wire g7760;
wire g4943;
wire g4587;
wire II12595;
wire g9260;
wire II12875;
wire g10795;
wire g6922;
wire g11580;
wire g5494;
wire g5215;
wire g8725;
wire g7028;
wire g6284;
wire II15568;
wire g6805;
wire g9884;
wire II12183;
wire g2522;
wire g7774;
wire g9702;
wire II14224;
wire g8070;
wire II17191;
wire g5756;
wire g2396;
wire II11261;
wire g7061;
wire g8404;
wire g6320;
wire g9729;
wire II10057;
wire g4620;
wire g9097;
wire II13212;
wire g10150;
wire g7889;
wire II8778;
wire g6404;
wire g10282;
wire g10119;
wire g7196;
wire g8841;
wire II9510;
wire g11276;
wire g8848;
wire g4986;
wire g8684;
wire g10580;
wire II12039;
wire g10034;
wire g9511;
wire g7278;
wire g3394;
wire g7907;
wire g8991;
wire g4398;
wire g2074;
wire g3810;
wire II14295;
wire g11596;
wire g6929;
wire g11313;
wire g11554;
wire g6202;
wire g4199;
wire II6517;
wire g4182;
wire II15959;
wire g11049;
wire g4069;
wire g2938;
wire g7675;
wire g9335;
wire g3281;
wire g4000;
wire g5194;
wire g8687;
wire g6819;
wire g6563;
wire II6761;
wire g4995;
wire g3062;
wire g8307;
wire g9389;
wire g6360;
wire II5751;
wire g10357;
wire II16514;
wire g5024;
wire g8968;
wire II7691;
wire g10179;
wire II14866;
wire g9900;
wire g7892;
wire II7684;
wire II10141;
wire g3774;
wire g9907;
wire g7089;
wire II4894;
wire II7683;
wire II14525;
wire g4355;
wire g7026;
wire g8447;
wire g4610;
wire g4940;
wire II7375;
wire g4396;
wire g6365;
wire g10195;
wire II12128;
wire g8191;
wire g7982;
wire g3412;
wire g10042;
wire II6501;
wire g8995;
wire II13300;
wire g3436;
wire II6331;
wire II7381;
wire II6827;
wire g6542;
wire g7763;
wire g9569;
wire II17347;
wire g10535;
wire g4556;
wire II10849;
wire g5729;
wire II5513;
wire II15400;
wire g2368;
wire g6561;
wire g4311;
wire g6293;
wire g5788;
wire g11249;
wire g11061;
wire g11238;
wire g6577;
wire g7911;
wire g6201;
wire II6106;
wire g5748;
wire g11305;
wire g5805;
wire g5216;
wire g11467;
wire g7352;
wire g11092;
wire g6629;
wire g5025;
wire II16607;
wire g7314;
wire g10913;
wire g2098;
wire II17202;
wire g10571;
wire g9785;
wire g2455;
wire g4342;
wire II17758;
wire g5445;
wire g4432;
wire g7367;
wire g3761;
wire g8361;
wire II7999;
wire g5680;
wire g4835;
wire g7030;
wire g4197;
wire g10666;
wire II13661;
wire II17121;
wire g6419;
wire g7696;
wire g8319;
wire g10561;
wire g11325;
wire g8892;
wire g6261;
wire II5722;
wire g8728;
wire g4009;
wire II14786;
wire g4236;
wire g2859;
wire g9715;
wire II11804;
wire g8532;
wire g10174;
wire g8403;
wire II6208;
wire II16571;
wire g3119;
wire g6872;
wire g2298;
wire g5498;
wire g5874;
wire g10550;
wire II5185;
wire g4401;
wire II9973;
wire g9879;
wire g7214;
wire g8119;
wire II5957;
wire g8170;
wire II12556;
wire II9673;
wire II14862;
wire II8529;
wire g7604;
wire g7073;
wire g11424;
wire g4454;
wire g3474;
wire g8780;
wire g10349;
wire g10417;
wire II12144;
wire g7192;
wire II16295;
wire g6853;
wire g8749;
wire g9594;
wire g7064;
wire g4212;
wire g4811;
wire g10176;
wire g8779;
wire II12907;
wire g7457;
wire g5983;
wire II15798;
wire g9849;
wire g8314;
wire g3067;
wire II7606;
wire II9769;
wire g4421;
wire g7895;
wire g6879;
wire II15205;
wire g6837;
wire g10681;
wire g3716;
wire g5743;
wire II7651;
wire g8075;
wire II15418;
wire g11437;
wire g7626;
wire g3404;
wire g6923;
wire II17704;
wire II6013;
wire g10784;
wire g5694;
wire g6994;
wire II11599;
wire II10974;
wire g7450;
wire g2018;
wire g9767;
wire g8385;
wire g6587;
wire g7938;
wire II16641;
wire g7523;
wire II15250;
wire II6941;
wire g6549;
wire II13515;
wire II10807;
wire g6523;
wire g4068;
wire II12199;
wire g4419;
wire g4526;
wire g4144;
wire g8757;
wire g4619;
wire g11595;
wire g8520;
wire II15956;
wire II8787;
wire II8358;
wire g4481;
wire g3333;
wire g4114;
wire g4756;
wire g6556;
wire g11514;
wire g3010;
wire II13200;
wire II14005;
wire g5758;
wire II8652;
wire g5478;
wire II5174;
wire g4839;
wire g4208;
wire g3438;
wire II10685;
wire g11034;
wire II5690;
wire g6951;
wire II14573;
wire g7936;
wire g10625;
wire II17719;
wire g2833;
wire II13027;
wire g6396;
wire g7991;
wire II17770;
wire g11507;
wire g9764;
wire II13194;
wire g2547;
wire II15033;
wire g6208;
wire g8787;
wire g7677;
wire g5814;
wire g10342;
wire II16387;
wire II16656;
wire g11009;
wire II7086;
wire II17505;
wire g7045;
wire II9221;
wire II11275;
wire g3399;
wire II5014;
wire g3768;
wire g7023;
wire II14873;
wire g11357;
wire II10322;
wire g3382;
wire g5541;
wire g5198;
wire g3912;
wire II10639;
wire II6360;
wire II9458;
wire g10374;
wire g8680;
wire g10366;
wire g9384;
wire g2356;
wire g5269;
wire g8766;
wire II16269;
wire g5629;
wire g9028;
wire g6055;
wire II16518;
wire g4266;
wire g2078;
wire g2915;
wire g9560;
wire g9750;
wire II7423;
wire II8388;
wire g4542;
wire g7539;
wire g10320;
wire g9317;
wire g8558;
wire g2112;
wire g4603;
wire g6093;
wire II16142;
wire g6185;
wire II15225;
wire g7219;
wire g1983;
wire II10355;
wire g4207;
wire II11814;
wire g8051;
wire g9951;
wire II13469;
wire g11401;
wire II14370;
wire g7925;
wire II14964;
wire g5047;
wire g10286;
wire II6792;
wire g3003;
wire g10254;
wire g5916;
wire g10471;
wire g11469;
wire g8186;
wire g2796;
wire g5536;
wire II11029;
wire g7321;
wire g2389;
wire II7889;
wire g5396;
wire g4803;
wire g7996;
wire II15608;
wire g3094;
wire g6239;
wire g4333;
wire g2534;
wire II17586;
wire II10240;
wire g3400;
wire II6965;
wire II5101;
wire g11540;
wire g11620;
wire g8324;
wire g9872;
wire g9515;
wire II17519;
wire II11647;
wire g4294;
wire g8045;
wire g7784;
wire g3077;
wire g9410;
wire II13442;
wire g8750;
wire g9361;
wire g3772;
wire II9380;
wire g2419;
wire II17724;
wire II15906;
wire II8543;
wire II6282;
wire g10499;
wire II10099;
wire g11168;
wire g11014;
wire g8004;
wire II12871;
wire g2450;
wire g2561;
wire II5166;
wire g3329;
wire g7680;
wire II13475;
wire g11558;
wire g8479;
wire II14914;
wire g4566;
wire II16720;
wire g11440;
wire g2847;
wire II12086;
wire II8797;
wire II15688;
wire g6857;
wire g7725;
wire g9935;
wire g11430;
wire g8033;
wire g6327;
wire g4880;
wire II10302;
wire II9062;
wire g5601;
wire g5548;
wire g10686;
wire g2719;
wire g9701;
wire g10523;
wire II14827;
wire g6434;
wire g4002;
wire g5527;
wire g10698;
wire II8606;
wire g9644;
wire g4012;
wire g8876;
wire g7202;
wire g9583;
wire II12469;
wire II6028;
wire II17216;
wire II13868;
wire g8064;
wire g2082;
wire g7379;
wire g10395;
wire g11649;
wire g5948;
wire g7817;
wire g2961;
wire II7408;
wire II16760;
wire II5529;
wire g8168;
wire g10578;
wire g11052;
wire II9836;
wire II10941;
wire g4387;
wire g10309;
wire g6301;
wire II16114;
wire g5996;
wire II12137;
wire g5191;
wire g6197;
wire g11389;
wire II12502;
wire II14194;
wire g9597;
wire g5203;
wire g11273;
wire II16897;
wire g4900;
wire g2980;
wire II5538;
wire g4259;
wire g7328;
wire g8302;
wire g11441;
wire g2248;
wire g4076;
wire g10726;
wire II6985;
wire g11419;
wire II6201;
wire g5177;
wire g7055;
wire g8246;
wire II15395;
wire g3506;
wire g5040;
wire g8716;
wire g10881;
wire g2515;
wire II11243;
wire g6226;
wire II13227;
wire g11310;
wire g8355;
wire g9808;
wire g5676;
wire II5378;
wire g4382;
wire II8738;
wire g11486;
wire g2850;
wire g9926;
wire II10374;
wire g10450;
wire g4225;
wire g4565;
wire g4188;
wire II12933;
wire g7052;
wire g7568;
wire II14697;
wire g8245;
wire g3661;
wire g5421;
wire g6420;
wire g7093;
wire II13639;
wire g4222;
wire II17675;
wire g5687;
wire g11609;
wire II12641;
wire g10231;
wire g2126;
wire g3829;
wire g4607;
wire II11829;
wire II7143;
wire II9282;
wire II17053;
wire g11185;
wire g10158;
wire g2116;
wire g9953;
wire II15756;
wire II16879;
wire g8068;
wire g6214;
wire g7821;
wire g10638;
wire II10623;
wire g6444;
wire II17610;
wire II7843;
wire g6355;
wire g7069;
wire g9261;
wire g9619;
wire g5004;
wire g5797;
wire g10474;
wire g2091;
wire g10731;
wire II7191;
wire II12076;
wire II11188;
wire g5085;
wire g10448;
wire g5515;
wire g4061;
wire II7735;
wire II10560;
wire g2343;
wire g8470;
wire g4096;
wire g5617;
wire II13295;
wire g9424;
wire II7112;
wire g8823;
wire g8970;
wire II15244;
wire g8412;
wire g11208;
wire II7321;
wire II10573;
wire II13460;
wire g3684;
wire II5815;
wire II13323;
wire g7905;
wire g10871;
wire II11263;
wire g4585;
wire g10467;
wire g3253;
wire g10878;
wire II13090;
wire g3290;
wire g2438;
wire g4502;
wire II12388;
wire g9708;
wire II8406;
wire II6196;
wire g6044;
wire g5846;
wire g9603;
wire II6468;
wire II17084;
wire II5809;
wire g6616;
wire g2906;
wire g11642;
wire II10831;
wire g2754;
wire g3782;
wire II17558;
wire II10508;
wire g2613;
wire II11071;
wire II12759;
wire II5684;
wire g5937;
wire g2243;
wire g4954;
wire II9953;
wire g10851;
wire II6226;
wire g9909;
wire g5492;
wire g11191;
wire II9174;
wire g6812;
wire II5254;
wire g2626;
wire g7635;
wire g9831;
wire g3106;
wire II12862;
wire g6102;
wire g9718;
wire g11471;
wire g4103;
wire g2179;
wire g9728;
wire II16413;
wire g6828;
wire g4723;
wire g10684;
wire g11231;
wire II9779;
wire g10518;
wire g2158;
wire II5383;
wire g11474;
wire g2104;
wire g11546;
wire II11767;
wire II12087;
wire g6817;
wire g8144;
wire g8516;
wire g4451;
wire g5499;
wire g5009;
wire g6535;
wire g7650;
wire g11016;
wire II10873;
wire g8972;
wire g2184;
wire g5319;
wire g9940;
wire g11111;
wire II12487;
wire g7943;
wire II10251;
wire II11904;
wire g6111;
wire g9447;
wire II12986;
wire g8646;
wire II6748;
wire g2800;
wire g4991;
wire g8507;
wire II9243;
wire II9829;
wire g4291;
wire g9354;
wire g10318;
wire g10929;
wire II7444;
wire g3743;
wire g4063;
wire g6135;
wire g6543;
wire g7562;
wire II15771;
wire II17633;
wire g7243;
wire g8118;
wire g7571;
wire g8703;
wire g4156;
wire g11643;
wire g4961;
wire II15548;
wire g9622;
wire g7556;
wire g11144;
wire g7804;
wire g2199;
wire II11159;
wire g11215;
wire g4479;
wire g8651;
wire g7606;
wire g3379;
wire g6427;
wire II5308;
wire II15458;
wire II8804;
wire g5914;
wire g6500;
wire g5250;
wire g6697;
wire gbuf4;
wire II9717;
wire II10584;
wire g9902;
wire g10482;
wire g10742;
wire g1993;
wire g5777;
wire g7508;
wire II9655;
wire g3220;
wire II17485;
wire II14340;
wire g6896;
wire II9402;
wire g5608;
wire g9474;
wire g10485;
wire II6546;
wire g8261;
wire II15804;
wire g8287;
wire g6271;
wire g6350;
wire g2844;
wire II5104;
wire II12913;
wire II16947;
wire g8642;
wire g8975;
wire g7757;
wire g9605;
wire g10753;
wire g8469;
wire g8462;
wire II7771;
wire II12251;
wire II6136;
wire g10311;
wire g9363;
wire g11343;
wire g8053;
wire II14270;
wire g4057;
wire g10133;
wire II11534;
wire g4898;
wire g7505;
wire g9869;
wire II12177;
wire II8780;
wire g8940;
wire g11031;
wire g9695;
wire II11701;
wire II7563;
wire II13648;
wire g4460;
wire II8561;
wire II17283;
wire g3696;
wire g7589;
wire g6268;
wire g10669;
wire g5936;
wire g10765;
wire g6663;
wire II13373;
wire II14349;
wire g4160;
wire g4932;
wire g4998;
wire II13412;
wire II5707;
wire II11312;
wire g7289;
wire g8239;
wire g8010;
wire g6125;
wire g6748;
wire g5006;
wire g2701;
wire g8164;
wire II15451;
wire g2839;
wire g9432;
wire II15323;
wire g5106;
wire II13747;
wire g2015;
wire II6870;
wire g4218;
wire g9610;
wire g8555;
wire II17374;
wire g4374;
wire g9573;
wire g8172;
wire II14185;
wire g8138;
wire g4675;
wire g11617;
wire g11634;
wire II9093;
wire g7290;
wire II9798;
wire g7536;
wire g11154;
wire g6738;
wire g2329;
wire g8884;
wire g4778;
wire II11037;
wire II15377;
wire II16867;
wire II16592;
wire II9156;
wire II10243;
wire g4865;
wire g6334;
wire g6755;
wire II9783;
wire g8383;
wire g11585;
wire g3683;
wire g9739;
wire g8437;
wire g10559;
wire g6744;
wire g7657;
wire g2550;
wire II6639;
wire g4716;
wire g6363;
wire g8025;
wire g5660;
wire g11339;
wire g8500;
wire g8105;
wire g10496;
wire g9240;
wire II8772;
wire II8795;
wire g9646;
wire II17470;
wire g7135;
wire II8664;
wire g6035;
wire II14543;
wire II5399;
wire g7595;
wire g10114;
wire g7298;
wire II5084;
wire II7648;
wire g5186;
wire g9680;
wire II9032;
wire g4884;
wire g10490;
wire g4126;
wire g7729;
wire II8996;
wire g8807;
wire g7131;
wire g7796;
wire g5981;
wire g1988;
wire g11574;
wire g2726;
wire g4966;
wire g10782;
wire II5451;
wire g2252;
wire g10334;
wire g5253;
wire g5943;
wire II12061;
wire g10923;
wire g6310;
wire II8839;
wire g9913;
wire g4414;
wire g9964;
wire II15586;
wire g7237;
wire g8736;
wire g6507;
wire II4917;
wire g10893;
wire II6664;
wire II14596;
wire g10793;
wire II5731;
wire g6156;
wire g6141;
wire II5501;
wire g7230;
wire g6236;
wire II13720;
wire II9409;
wire g11492;
wire g7615;
wire g8663;
wire g2882;
wire g7592;
wire II6166;
wire g3704;
wire II14681;
wire g7662;
wire II10461;
wire II16079;
wire g4047;
wire g9125;
wire II14352;
wire g2372;
wire g4733;
wire g6219;
wire II13114;
wire g7669;
wire g11456;
wire II6513;
wire II6802;
wire II10655;
wire g2202;
wire II11964;
wire II15335;
wire g4821;
wire g10504;
wire g5863;
wire g11088;
wire g6417;
wire g7971;
wire g3326;
wire g2335;
wire II10054;
wire g7148;
wire g8630;
wire II11740;
wire II5737;
wire g6144;
wire g4682;
wire g7786;
wire II8670;
wire II13794;
wire g2042;
wire g8036;
wire II12021;
wire g10164;
wire g10383;
wire II17164;
wire II15045;
wire II15999;
wire g6464;
wire g10546;
wire g6572;
wire g7477;
wire II6159;
wire g9009;
wire II15293;
wire g10278;
wire g8277;
wire g5485;
wire g7913;
wire g10717;
wire g2212;
wire II7920;
wire g6048;
wire g5531;
wire g2223;
wire g4670;
wire g7144;
wire II9688;
wire g8294;
wire II16487;
wire II5629;
wire II12366;
wire g6883;
wire g10544;
wire II11974;
wire II9338;
wire g8890;
wire g5035;
wire II11296;
wire g6803;
wire g11021;
wire II6979;
wire g11614;
wire g11172;
wire g8399;
wire g7441;
wire g5524;
wire g10223;
wire II8728;
wire II16363;
wire g11350;
wire g8198;
wire g11551;
wire g10528;
wire g8425;
wire II13776;
wire g9686;
wire II7048;
wire g8925;
wire g10197;
wire II6495;
wire II10445;
wire II12644;
wire g7682;
wire g6655;
wire g10864;
wire II6264;
wire g6710;
wire g8363;
wire g9824;
wire g7850;
wire g8845;
wire g7008;
wire II9558;
wire II9605;
wire g6117;
wire II13859;
wire g5166;
wire g7388;
wire II12229;
wire g2024;
wire g11219;
wire II7417;
wire g4636;
wire g7733;
wire g11345;
wire II12765;
wire II5282;
wire g10751;
wire g10971;
wire g7882;
wire g8667;
wire g6175;
wire g8616;
wire g11483;
wire II5728;
wire g5821;
wire g5143;
wire g6930;
wire g5211;
wire g3052;
wire II10274;
wire II6911;
wire II15214;
wire II5926;
wire g10763;
wire II17312;
wire g7317;
wire II10282;
wire II17306;
wire II11383;
wire II12457;
wire g5196;
wire g7385;
wire g6085;
wire g4467;
wire g6720;
wire II16000;
wire II8379;
wire g9452;
wire g10758;
wire g4805;
wire g2273;
wire II11394;
wire g8767;
wire II14906;
wire g6554;
wire g7849;
wire g5245;
wire II13314;
wire g2917;
wire g6450;
wire g11240;
wire II11241;
wire g110;
wire II6487;
wire g2038;
wire II13376;
wire II13273;
wire g9947;
wire g5218;
wire g6915;
wire g3301;
wire g4769;
wire II14876;
wire II14694;
wire II7269;
wire g7432;
wire g10948;
wire g7331;
wire II12376;
wire g10771;
wire II15257;
wire g3946;
wire g8132;
wire g5075;
wire g3161;
wire II4866;
wire II16007;
wire g4189;
wire g7357;
wire II7876;
wire g7965;
wire g10126;
wire g4093;
wire g7188;
wire II9046;
wire gbuf2;
wire g9531;
wire II13553;
wire II10102;
wire g9835;
wire g10508;
wire II15162;
wire II11614;
wire g2407;
wire g5883;
wire g6701;
wire II7035;
wire II8285;
wire g11079;
wire g10264;
wire II6324;
wire g10779;
wire g8622;
wire II7411;
wire g1990;
wire II5050;
wire g4789;
wire g2646;
wire II5469;
wire g7306;
wire g8151;
wire g2579;
wire g2174;
wire g2542;
wire g10454;
wire II15266;
wire II13259;
wire g7342;
wire g3729;
wire g7269;
wire II9096;
wire g4436;
wire g4509;
wire II14579;
wire g5623;
wire g10462;
wire g11300;
wire II13209;
wire II11318;
wire II11845;
wire II13309;
wire g11195;
wire II17368;
wire g10062;
wire g11109;
wire g3992;
wire g7746;
wire II12442;
wire g3374;
wire g9928;
wire g4443;
wire g3629;
wire II6716;
wire II8161;
wire g4429;
wire g10723;
wire II13249;
wire g8814;
wire II13785;
wire g5725;
wire g11296;
wire II9168;
wire g10537;
wire g11285;
wire g10141;
wire g3586;
wire g11221;
wire II6569;
wire II5932;
wire II13089;
wire g3089;
wire g10091;
wire g6622;
wire g6109;
wire g10652;
wire II11926;
wire g4472;
wire II12490;
wire II11698;
wire g6319;
wire II16856;
wire II7459;
wire g3720;
wire g11162;
wire II11303;
wire II17142;
wire II7523;
wire II5289;
wire g9877;
wire II9256;
wire g10153;
wire g9599;
wire g5595;
wire g8782;
wire g3143;
wire g10530;
wire g9344;
wire II5986;
wire g3516;
wire g3458;
wire g10148;
wire g4053;
wire II9483;
wire II8626;
wire II6309;
wire II12296;
wire g4975;
wire II8903;
wire g8921;
wire g11422;
wire g6940;
wire II5077;
wire II16723;
wire II8410;
wire g10912;
wire g4712;
wire g4758;
wire II8650;
wire g11612;
wire II15514;
wire g3583;
wire g6568;
wire g10582;
wire g6063;
wire g8695;
wire g7975;
wire II9253;
wire g6529;
wire g3529;
wire g6191;
wire g10908;
wire g5276;
wire II11225;
wire II7205;
wire g5992;
wire g4363;
wire g10557;
wire g8077;
wire g10376;
wire g9417;
wire g11093;
wire II14564;
wire g6454;
wire II16953;
wire II12168;
wire II9591;
wire g7781;
wire g8954;
wire g4412;
wire g11247;
wire g7768;
wire g5068;
wire g5752;
wire g6431;
wire g8226;
wire II4995;
wire g6300;
wire g11512;
wire II9440;
wire II6256;
wire II13577;
wire II17642;
wire g8096;
wire II15380;
wire g5994;
wire II13385;
wire g2524;
wire g10456;
wire g4238;
wire II7220;
wire II8724;
wire II10162;
wire g8882;
wire g4417;
wire II12196;
wire g5696;
wire g10353;
wire g10137;
wire g9151;
wire g6558;
wire g9673;
wire g1999;
wire II5740;
wire II8751;
wire II12849;
wire g10905;
wire g5823;
wire II5576;
wire II15488;
wire II12123;
wire II12279;
wire II17669;
wire II11996;
wire g9386;
wire II5358;
wire g2549;
wire g6398;
wire II15908;
wire g8357;
wire g3354;
wire g6534;
wire II16647;
wire g4066;
wire g5230;
wire II10278;
wire g8139;
wire II6260;
wire g4583;
wire II7399;
wire g6589;
wire g4772;
wire II9383;
wire II15235;
wire II16784;
wire g10593;
wire g4631;
wire II10075;
wire II11076;
wire II9762;
wire g7078;
wire g3820;
wire g8789;
wire g7903;
wire g7043;
wire II5149;
wire g5476;
wire g10747;
wire II6891;
wire II13360;
wire g7146;
wire g5850;
wire II5611;
wire II9208;
wire II9087;
wire II5843;
wire g4366;
wire g7096;
wire g7989;
wire g10364;
wire g7679;
wire g2016;
wire g7347;
wire II11326;
wire II13627;
wire g6183;
wire g9736;
wire II15855;
wire II17350;
wire g11047;
wire g8541;
wire g9527;
wire g8445;
wire g7010;
wire g9509;
wire II17100;
wire g4109;
wire g4394;
wire II11135;
wire II13005;
wire g10304;
wire g5681;
wire g10858;
wire g3275;
wire II14690;
wire II6337;
wire II9567;
wire g6684;
wire g11332;
wire II13020;
wire II17537;
wire II13522;
wire g11583;
wire II17636;
wire gbuf9;
wire g4292;
wire II9479;
wire g7312;
wire g9866;
wire g11214;
wire g10627;
wire II6794;
wire II5348;
wire II9006;
wire II6177;
wire II9013;
wire g7609;
wire II16087;
wire g3268;
wire g7778;
wire II6836;
wire II11055;
wire II13105;
wire g3364;
wire II17701;
wire II5850;
wire g5546;
wire g6878;
wire g5309;
wire II9053;
wire II6338;
wire II16149;
wire g7365;
wire II17182;
wire II5518;
wire g7801;
wire II7154;
wire g5513;
wire II13293;
wire g5733;
wire g11454;
wire g5767;
wire g4378;
wire II7366;
wire II5351;
wire g4340;
wire g9889;
wire g10193;
wire g6281;
wire g10888;
wire g7138;
wire g5418;
wire g8309;
wire g10361;
wire II12776;
wire g2351;
wire g8428;
wire g11593;
wire g11270;
wire II10153;
wire II17228;
wire g11005;
wire II17288;
wire II7342;
wire g2228;
wire g10761;
wire II8456;
wire g3186;
wire II9684;
wire g10122;
wire II16330;
wire g9820;
wire g3532;
wire g4186;
wire g10189;
wire g2119;
wire g4314;
wire g3983;
wire g2798;
wire g4329;
wire g9933;
wire II17194;
wire II11756;
wire g9263;
wire g7897;
wire g4958;
wire g7212;
wire g3414;
wire g4837;
wire II6273;
wire g10172;
wire II16261;
wire II15523;
wire II5862;
wire II4956;
wire g4992;
wire II15329;
wire g3406;
wire g7359;
wire g2853;
wire g4004;
wire II10651;
wire II13828;
wire II8715;
wire g8401;
wire g8874;
wire g7602;
wire II6409;
wire g11071;
wire g2752;
wire g7190;
wire II16531;
wire g6815;
wire g6198;
wire II17258;
wire II9625;
wire g9339;
wire g7062;
wire II14948;
wire g10031;
wire II12094;
wire g9713;
wire g6830;
wire g8777;
wire g10805;
wire g4380;
wire g8747;
wire g10144;
wire g6839;
wire g6228;
wire g9955;
wire g5649;
wire II7255;
wire g2802;
wire g8248;
wire g4551;
wire g8821;
wire g8826;
wire g4220;
wire g3663;
wire II10610;
wire g5857;
wire g4488;
wire g8523;
wire g8802;
wire g10740;
wire II15503;
wire II14202;
wire g11181;
wire g2421;
wire II8133;
wire g7197;
wire g10869;
wire II11873;
wire g2118;
wire II15601;
wire g4951;
wire g4456;
wire g7670;
wire II12363;
wire g11058;
wire II8007;
wire II11722;
wire II11433;
wire II6125;
wire g2791;
wire II8098;
wire g7426;
wire g8376;
wire II5973;
wire g5741;
wire II11194;
wire II13744;
wire g10786;
wire g7808;
wire g10182;
wire II11180;
wire g10437;
wire g11626;
wire g8670;
wire g8718;
wire II7104;
wire g7825;
wire g6913;
wire II9120;
wire g2268;
wire g2432;
wire II12598;
wire g4257;
wire II14400;
wire g2439;
wire g10724;
wire II12215;
wire g10275;
wire g11488;
wire II13816;
wire g9310;
wire g11601;
wire g9895;
wire II17051;
wire g4371;
wire g10414;
wire II7865;
wire g4227;
wire g4327;
wire g9906;
wire II13122;
wire g4536;
wire g5391;
wire II10769;
wire g5128;
wire g4749;
wire II14211;
wire g6618;
wire g4335;
wire II7450;
wire g9091;
wire II16534;
wire II5258;
wire g8945;
wire g4195;
wire g8764;
wire II13077;
wire g2275;
wire g6729;
wire g7354;
wire g5910;
wire g8240;
wire g9422;
wire g2818;
wire II8199;
wire II4873;
wire g6321;
wire g2813;
wire g5233;
wire g5222;
wire g3273;
wire II10771;
wire g6206;
wire g10428;
wire II15986;
wire II12004;
wire g8449;
wire II11289;
wire II15284;
wire II16370;
wire g7546;
wire II12910;
wire g3522;
wire II13099;
wire II13902;
wire II7662;
wire g7001;
wire g10050;
wire g5001;
wire g5171;
wire II13894;
wire II11357;
wire g3989;
wire g9108;
wire g7633;
wire g3434;
wire g2908;
wire g3256;
wire g3710;
wire II8762;
wire II12829;
wire II6421;
wire g8797;
wire g10263;
wire g5703;
wire II17695;
wire g7067;
wire g8639;
wire g4006;
wire g8066;
wire II16769;
wire II6436;
wire g8576;
wire g5642;
wire g2892;
wire g5848;
wire g7815;
wire g2096;
wire g11628;
wire II7713;
wire g2743;
wire II15708;
wire g10252;
wire g10281;
wire g2166;
wire g4430;
wire II14552;
wire II13185;
wire g8783;
wire g11656;
wire g1981;
wire g8047;
wire g2073;
wire g7628;
wire II17487;
wire II8192;
wire II17268;
wire g6313;
wire g8711;
wire II17295;
wire g5836;
wire g11445;
wire II5323;
wire II16059;
wire II6553;
wire g4763;
wire II17321;
wire g10203;
wire II17681;
wire II17401;
wire g4500;
wire g8628;
wire g9859;
wire g6956;
wire g7224;
wire g11407;
wire II14303;
wire g9870;
wire g7753;
wire II11508;
wire II11501;
wire g6751;
wire g6240;
wire II16379;
wire g10297;
wire g5529;
wire II9662;
wire II17188;
wire g6693;
wire II12003;
wire g9651;
wire II9248;
wire g3261;
wire II7185;
wire g8598;
wire g8415;
wire g4609;
wire g8162;
wire II13329;
wire g3815;
wire II6576;
wire g10307;
wire g2555;
wire g6842;
wire II7233;
wire g8602;
wire g10430;
wire g4205;
wire II13367;
wire II10813;
wire g4561;
wire g6514;
wire g5201;
wire g6151;
wire g4558;
wire g3756;
wire g6361;
wire g11103;
wire II7276;
wire II10901;
wire g6644;
wire II10394;
wire g7200;
wire g7071;
wire g2001;
wire g4949;
wire g10393;
wire II13347;
wire g11387;
wire g8342;
wire g9775;
wire II12655;
wire II8985;
wire g6705;
wire g7998;
wire g5193;
wire g1973;
wire g10347;
wire g8790;
wire g2084;
wire g4783;
wire g11390;
wire II13338;
wire g2777;
wire g5575;
wire II9810;
wire g10521;
wire g4492;
wire II12517;
wire g6014;
wire g5892;
wire g2296;
wire II5341;
wire g4306;
wire II14140;
wire II13513;
wire II13388;
wire g7723;
wire II8604;
wire g7327;
wire g4575;
wire II7213;
wire g9649;
wire II9368;
wire g7039;
wire g4889;
wire g11050;
wire g4512;
wire g8175;
wire II10719;
wire g10576;
wire II8293;
wire II13878;
wire g6715;
wire g7205;
wire g9841;
wire II14277;
wire II13166;
wire II17413;
wire g5052;
wire g4010;
wire II8204;
wire g4896;
wire g8510;
wire II9901;
wire g5612;
wire g5444;
wire g2013;
wire II9930;
wire g10250;
wire II16811;
wire g5148;
wire g7587;
wire g4874;
wire g7520;
wire g9585;
wire II12571;
wire g5280;
wire II5279;
wire g5179;
wire g6299;
wire II7249;
wire II13711;
wire g8800;
wire g10464;
wire II6666;
wire II12403;
wire g10408;
wire g2593;
wire g8677;
wire g3212;
wire II10072;
wire g11299;
wire II10381;
wire g6258;
wire g10895;
wire g8427;
wire g3215;
wire II15171;
wire II12484;
wire II11173;
wire II17510;
wire g5737;
wire g5812;
wire II7447;
wire g3208;
wire g6262;
wire g4882;
wire g3681;
wire g6231;
wire II17742;
wire g3914;
wire II10221;
wire g2330;
wire g6123;
wire II5245;
wire g6592;
wire g10494;
wire g6336;
wire g6171;
wire g8213;
wire II5497;
wire g7534;
wire g10233;
wire g7263;
wire g10268;
wire g6798;
wire II16046;
wire II11731;
wire II17749;
wire g8965;
wire g9915;
wire g9367;
wire II9265;
wire II10138;
wire g11632;
wire g10791;
wire g6901;
wire g2728;
wire g2057;
wire II10084;
wire g3105;
wire II9801;
wire II12012;
wire g2086;
wire g5050;
wire g11038;
wire g5184;
wire g5794;
wire g9290;
wire g3861;
wire g11538;
wire g11509;
wire g7296;
wire g4128;
wire g3939;
wire g8699;
wire g6746;
wire II4980;
wire g2981;
wire g5304;
wire II14802;
wire II10526;
wire g10214;
wire g4117;
wire g6107;
wire g8381;
wire g8023;
wire g2775;
wire g8486;
wire II17466;
wire II9185;
wire g11500;
wire g7794;
wire g7235;
wire g6158;
wire g9737;
wire g11160;
wire g9843;
wire g4759;
wire II17569;
wire g4714;
wire g6330;
wire II9727;
wire II13765;
wire g6295;
wire g2650;
wire g8124;
wire g4677;
wire g6974;
wire g9273;
wire g3384;
wire II8820;
wire g7664;
wire II8563;
wire g11267;
wire g8055;
wire II16598;
wire g4169;
wire g6312;
wire II13735;
wire II6046;
wire II10174;
wire g9980;
wire g8280;
wire II8740;
wire g9863;
wire g10135;
wire g11330;
wire II13915;
wire g10238;
wire g4059;
wire g4752;
wire g8937;
wire II16982;
wire g2695;
wire g8019;
wire g11572;
wire II15580;
wire g4277;
wire II14490;
wire g10295;
wire g4548;
wire II16475;
wire g2320;
wire II12258;
wire g8756;
wire g3630;
wire g2003;
wire II9720;
wire g8107;
wire II11097;
wire g9777;
wire II13260;
wire II12068;
wire II10180;
wire II5638;
wire II11367;
wire g10708;
wire g5656;
wire g5667;
wire g6892;
wire II14751;
wire g3770;
wire g5102;
wire g8142;
wire g11461;
wire g8000;
wire g5265;
wire g7613;
wire II5023;
wire g9705;
wire II15820;
wire g7338;
wire II5316;
wire II11068;
wire g11233;
wire g3512;
wire g2496;
wire g7241;
wire II8892;
wire g10502;
wire II15725;
wire II9068;
wire g9904;
wire II5719;
wire II5057;
wire g3539;
wire g4386;
wire g5292;
wire g2178;
wire g6115;
wire II6363;
wire II8842;
wire II10234;
wire II12817;
wire g4477;
wire g4373;
wire II12796;
wire g4552;
wire II17161;
wire g11017;
wire g7427;
wire g9833;
wire g2955;
wire II11387;
wire g5724;
wire g4736;
wire II13280;
wire II9749;
wire g6795;
wire g11257;
wire II12107;
wire g7879;
wire g8517;
wire II5449;
wire g6277;
wire II10126;
wire g11010;
wire II12047;
wire II6523;
wire II6168;
wire g7410;
wire II11494;
wire II4900;
wire II5092;
wire II13857;
wire g2944;
wire g10259;
wire g10738;
wire II6449;
wire g11645;
wire g6100;
wire g10329;
wire g6810;
wire g2410;
wire g5518;
wire g4337;
wire II11683;
wire II6351;
wire g5773;
wire g2105;
wire II15453;
wire g8122;
wire g8129;
wire II15826;
wire g6110;
wire g6993;
wire g8509;
wire g6352;
wire II10930;
wire g10927;
wire g2172;
wire g2689;
wire II12712;
wire g3390;
wire II9452;
wire g11271;
wire g8644;
wire II10087;
wire II14412;
wire II4930;
wire g9624;
wire II13945;
wire II15872;
wire g8943;
wire g5226;
wire g6506;
wire g11410;
wire g7847;
wire II13621;
wire g7712;
wire g4211;
wire g2156;
wire g3369;
wire II8929;
wire II5798;
wire g6699;
wire II11759;
wire II5486;
wire g9837;
wire g8931;
wire g4158;
wire g7284;
wire II11914;
wire II5946;
wire g10155;
wire II9536;
wire g4080;
wire II16015;
wire II10914;
wire g9420;
wire g2271;
wire g9272;
wire g6181;
wire g7304;
wire g4308;
wire II15392;
wire g5638;
wire g3750;
wire g7186;
wire II6417;
wire II7014;
wire g6925;
wire g2123;
wire II17394;
wire g6446;
wire g10662;
wire II11510;
wire g4445;
wire g10849;
wire g2207;
wire g9328;
wire g11040;
wire g1968;
wire g10510;
wire II15247;
wire g5533;
wire II10063;
wire g5604;
wire II13660;
wire g8332;
wire II12607;
wire II9866;
wire II10864;
wire g6075;
wire II7323;
wire g2867;
wire g3336;
wire II10852;
wire II6856;
wire II6999;
wire g6730;
wire g6307;
wire g7963;
wire g5881;
wire g8796;
wire g9946;
wire g5895;
wire g11068;
wire II16635;
wire g2445;
wire g3497;
wire g6253;
wire II5292;
wire g3904;
wire II11299;
wire II16688;
wire II14264;
wire g8304;
wire II13552;
wire g9612;
wire g5108;
wire g11615;
wire g4915;
wire g2190;
wire g7511;
wire g10721;
wire II16616;
wire II5020;
wire II6489;
wire g2889;
wire g10506;
wire g2827;
wire g8431;
wire g5011;
wire g6821;
wire g11007;
wire g4679;
wire II8126;
wire II6474;
wire g11298;
wire g8648;
wire g8134;
wire II12475;
wire g3784;
wire II13302;
wire II16067;
wire g3734;
wire g3141;
wire II5371;
wire g6876;
wire g6742;
wire g5889;
wire II11581;
wire g4364;
wire g5345;
wire II13717;
wire g4427;
wire II10499;
wire g6898;
wire g6441;
wire g6481;
wire g9875;
wire II11065;
wire g9392;
wire II5675;
wire g10044;
wire g5662;
wire g6703;
wire II11423;
wire II12853;
wire g4470;
wire g4973;
wire g11077;
wire g2254;
wire g6620;
wire II17492;
wire g11499;
wire II13546;
wire g3732;
wire g3944;
wire g7454;
wire II14097;
wire g8951;
wire g7951;
wire g5259;
wire g2855;
wire II9642;
wire g4264;
wire II11408;
wire g11193;
wire g4779;
wire II6299;
wire g4507;
wire II6507;
wire g2214;
wire g7941;
wire II13036;
wire g10853;
wire g9419;
wire g8654;
wire g6885;
wire g5066;
wire g10166;
wire g6405;
wire g5746;
wire g11544;
wire g2884;
wire g10001;
wire g7885;
wire II17460;
wire g10598;
wire II10484;
wire g6634;
wire II9293;
wire II11833;
wire II12562;
wire g7142;
wire g2050;
wire g2221;
wire g4731;
wire g10385;
wire II11531;
wire g2044;
wire II15424;
wire II9080;
wire II12948;
wire g6083;
wire II11659;
wire g6346;
wire II17549;
wire g4616;
wire II8480;
wire II13797;
wire g10548;
wire II17096;
wire g2241;
wire g5504;
wire g4725;
wire II11127;
wire g7102;
wire II8328;
wire g5627;
wire g3584;
wire II4997;
wire II16763;
wire II11947;
wire II7749;
wire g8923;
wire II17459;
wire g7766;
wire g6286;
wire g7048;
wire II7033;
wire g10107;
wire g8502;
wire g11170;
wire g5030;
wire II10334;
wire g7984;
wire g11402;
wire II11235;
wire g5261;
wire g2204;
wire g7755;
wire g10331;
wire II16098;
wire II15768;
wire g6656;
wire g3417;
wire g8380;
wire g10866;
wire g10777;
wire g4282;
wire g10604;
wire g9740;
wire g4194;
wire g4510;
wire g4823;
wire g5865;
wire II6879;
wire II5007;
wire II5395;
wire g7363;
wire II17522;
wire g7731;
wire g7956;
wire g4140;
wire g9807;
wire g11020;
wire g5111;
wire g8582;
wire g11369;
wire g3092;
wire g3335;
wire II14312;
wire II15598;
wire g6224;
wire g6980;
wire g10526;
wire g4284;
wire II8835;
wire II14379;
wire g7460;
wire g5819;
wire II9854;
wire II6322;
wire g6462;
wire II10716;
wire g8059;
wire II16469;
wire g7439;
wire II11783;
wire g2068;
wire g8660;
wire g7467;
wire II7674;
wire g5098;
wire g3875;
wire g11360;
wire II10601;
wire g3352;
wire II10713;
wire g7345;
wire II17296;
wire II8215;
wire g8255;
wire g8365;
wire g6082;
wire II15464;
wire II10340;
wire g6672;
wire g11261;
wire II13674;
wire g6089;
wire g6967;
wire g9030;
wire g6777;
wire g5037;
wire II12303;
wire g7915;
wire II6034;
wire II9896;
wire g7472;
wire g8224;
wire II8934;
wire II12835;
wire g7708;
wire g2950;
wire g6960;
wire g11095;
wire g2759;
wire g4738;
wire g8611;
wire g4338;
wire g3706;
wire II9029;
wire g11327;
wire g8196;
wire II13433;
wire g3759;
wire g10370;
wire g11639;
wire g10355;
wire g9343;
wire II7654;
wire g2374;
wire II7099;
wire g7684;
wire g3056;
wire g7020;
wire II12586;
wire g2444;
wire g7288;
wire g8063;
wire g9414;
wire g10807;
wire II13708;
wire g10226;
wire II13779;
wire g11508;
wire g2095;
wire II6838;
wire g8273;
wire g7509;
wire II4859;
wire II8403;
wire g4324;
wire g3322;
wire g6712;
wire II11989;
wire II12978;
wire II6757;
wire g2185;
wire g9829;
wire g6686;
wire II11710;
wire II14982;
wire g6471;
wire g11334;
wire II9848;
wire g8253;
wire II5919;
wire g11381;
wire g4397;
wire II15386;
wire g2920;
wire II17567;
wire II8803;
wire II11444;
wire g9529;
wire g10868;
wire II6770;
wire g7360;
wire g8049;
wire g4944;
wire g7614;
wire g8849;
wire g3047;
wire g1987;
wire II11342;
wire g7277;
wire g8610;
wire g2997;
wire II15604;
wire II17297;
wire gbuf12;
wire g7037;
wire g5110;
wire g3395;
wire II13409;
wire g6825;
wire g7226;
wire g10013;
wire g9076;
wire II9514;
wire II4777;
wire g10324;
wire g2434;
wire II7453;
wire g6788;
wire g2237;
wire II14888;
wire g5838;
wire g7887;
wire g3423;
wire II7173;
wire II9129;
wire II8591;
wire g6522;
wire g9391;
wire g11184;
wire g3371;
wire g9679;
wire g8872;
wire g5593;
wire II16735;
wire g11396;
wire g4904;
wire II14612;
wire II12002;
wire g6305;
wire II16072;
wire g4051;
wire II16492;
wire g3980;
wire g5173;
wire g4104;
wire g5736;
wire II17692;
wire g9556;
wire g10391;
wire II12505;
wire g6869;
wire g7728;
wire g8889;
wire g10351;
wire g8869;
wire g9607;
wire II8605;
wire g4202;
wire g6516;
wire g11405;
wire g8009;
wire g10064;
wire g7721;
wire II13636;
wire g8235;
wire g9892;
wire II13043;
wire g4464;
wire g4907;
wire II17450;
wire II6288;
wire g4229;
wire g5858;
wire g3008;
wire II6110;
wire II14279;
wire g2261;
wire II14540;
wire g11490;
wire II11008;
wire g6221;
wire g6424;
wire g6680;
wire II16252;
wire g6386;
wire g7672;
wire g10629;
wire g9857;
wire g4994;
wire II13102;
wire g5644;
wire g8724;
wire g5264;
wire g9352;
wire II7345;
wire g8344;
wire g6242;
wire g5122;
wire II16273;
wire g11056;
wire g10423;
wire II8340;
wire II5960;
wire II9669;
wire II11921;
wire II6989;
wire g5503;
wire g6068;
wire II4961;
wire g6449;
wire II5264;
wire g5762;
wire g9590;
wire g9896;
wire g8156;
wire g6440;
wire II5821;
wire g10800;
wire II13250;
wire g5678;
wire g2233;
wire g10553;
wire II10388;
wire g6933;
wire II6851;
wire g7270;
wire g8824;
wire g7341;
wire II10195;
wire g7203;
wire II12009;
wire g4254;
wire g10584;
wire II7817;
wire g2793;
wire II12529;
wire II7315;
wire II7829;
wire g6187;
wire II15196;
wire g7718;
wire g9965;
wire II7847;
wire II11626;
wire II15635;
wire g5661;
wire g8607;
wire g9958;
wire g11158;
wire II7625;
wire g5801;
wire g6574;
wire II12971;
wire II16080;
wire g4299;
wire g8952;
wire II14918;
wire II9737;
wire II14306;
wire II11728;
wire g8475;
wire g10634;
wire II12075;
wire II16175;
wire II12133;
wire II13901;
wire g6040;
wire II6754;
wire II14136;
wire g6311;
wire II12751;
wire II5271;
wire g11624;
wire g11448;
wire II10305;
wire g7403;
wire g4322;
wire g4877;
wire II6590;
wire II12029;
wire II15241;
wire g2122;
wire g7419;
wire II10753;
wire g5044;
wire g4953;
wire g9106;
wire g7376;
wire g9850;
wire g5220;
wire II12081;
wire g8721;
wire II16808;
wire II10027;
wire g5511;
wire II9202;
wire g11180;
wire II5036;
wire g6438;
wire g11289;
wire II14045;
wire g7126;
wire II16742;
wire g8592;
wire g8579;
wire g7742;
wire g8793;
wire g8574;
wire g6210;
wire g7324;
wire g5392;
wire g2511;
wire g2499;
wire II17281;
wire g10298;
wire g2518;
wire g8438;
wire g9804;
wire g4719;
wire g10479;
wire II17344;
wire g7420;
wire II11817;
wire g6342;
wire g5090;
wire g11204;
wire g9554;
wire g9409;
wire g8442;
wire II10733;
wire g2909;
wire g11373;
wire g11434;
wire II6055;
wire II9461;
wire g7098;
wire II15344;
wire g6165;
wire g6911;
wire II12520;
wire g7583;
wire II17112;
wire g9616;
wire g7210;
wire g10809;
wire g6265;
wire g2075;
wire II9677;
wire g8174;
wire II10996;
wire g7899;
wire II12108;
wire g8969;
wire g2820;
wire II7593;
wire g5654;
wire g6359;
wire g5722;
wire II13224;
wire g4588;
wire g7336;
wire II11797;
wire II14989;
wire II6762;
wire g9781;
wire II7357;
wire II8308;
wire II12339;
wire g7218;
wire g10191;
wire g7348;
wire g10711;
wire g8785;
wire II6102;
wire II16787;
wire II16805;
wire II10159;
wire g5878;
wire g11352;
wire II7996;
wire II13586;
wire II12538;
wire g3981;
wire g10903;
wire g11255;
wire II14958;
wire II9305;
wire g8775;
wire g3284;
wire g6625;
wire g3330;
wire g8604;
wire g8713;
wire II17493;
wire g10302;
wire g8760;
wire g3266;
wire II10060;
wire II16373;
wire II7793;
wire g2108;
wire g5759;
wire g5740;
wire g11606;
wire g2843;
wire g6954;
wire g6840;
wire g8110;
wire g8417;
wire g6862;
wire II8752;
wire g11189;
wire g4183;
wire g6566;
wire g8688;
wire g2399;
wire g9882;
wire II15814;
wire g5095;
wire II17773;
wire g8306;
wire g9712;
wire g7901;
wire g4346;
wire g2902;
wire g2226;
wire g2958;
wire g10291;
wire II15036;
wire g8407;
wire g11588;
wire II13400;
wire g4834;
wire II6777;
wire g3906;
wire II11770;
wire g11201;
wire II10979;
wire g2364;
wire II15353;
wire g10821;
wire g11210;
wire g11319;
wire g2382;
wire II7336;
wire g9772;
wire g10288;
wire II11593;
wire g2390;
wire g9704;
wire II15763;
wire II17393;
wire g6128;
wire g6283;
wire II16184;
wire g8366;
wire g3416;
wire g8056;
wire II12120;
wire g3353;
wire II17252;
wire g4216;
wire g6640;
wire II15592;
wire g3530;
wire g3479;
wire g10663;
wire g8772;
wire gbuf7;
wire II10822;
wire g6794;
wire II7369;
wire g6052;
wire g11590;
wire g9822;
wire g3811;
wire II7852;
wire g5697;
wire g11149;
wire g7060;
wire g11392;
wire g8957;
wire g9763;
wire g10928;
wire g4525;
wire g2883;
wire g10460;
wire g4987;
wire g11277;
wire g2004;
wire II9349;
wire g8378;
wire g4638;
wire II6498;
wire g6527;
wire g7891;
wire g11245;
wire II11115;
wire g8071;
wire g3386;
wire g8842;
wire g10033;
wire II5992;
wire g7992;
wire II7909;
wire g7806;
wire II13867;
wire g3693;
wire II5053;
wire II5916;
wire g6091;
wire g8990;
wire g11597;
wire g4640;
wire II9056;
wire g11101;
wire g11037;
wire g3362;
wire II12547;
wire g11314;
wire II9822;
wire g6205;
wire II11279;
wire g2454;
wire g2459;
wire g7621;
wire II14509;
wire g9506;
wire g6778;
wire g11217;
wire II11719;
wire g6289;
wire g9908;
wire g6895;
wire g7813;
wire II11467;
wire g4232;
wire II6686;
wire g6583;
wire g9931;
wire II11217;
wire g6591;
wire g6182;
wire II10165;
wire g11503;
wire II8031;
wire II12326;
wire II13812;
wire g7977;
wire II5935;
wire II7295;
wire II8730;
wire II7006;
wire II6480;
wire g7195;
wire g9664;
wire g3775;
wire g8317;
wire II14182;
wire g5980;
wire g8040;
wire II13109;
wire g10346;
wire II5203;
wire II8039;
wire g7356;
wire g11328;
wire g9692;
wire g3763;
wire II7378;
wire g2303;
wire g7608;
wire g7041;
wire g7526;
wire g6059;
wire II13290;
wire g9349;
wire g10449;
wire g10205;
wire g7932;
wire g11078;
wire g4362;
wire II15302;
wire II15479;
wire g9732;
wire II9371;
wire g10621;
wire II9043;
wire g11269;
wire g6763;
wire g7987;
wire g10802;
wire g4604;
wire g8116;
wire g10442;
wire II7291;
wire g10489;
wire g7042;
wire II11587;
wire g3432;
wire g6132;
wire g5474;
wire g9760;
wire II5940;
wire g4008;
wire g5852;
wire g9860;
wire II11091;
wire g5754;
wire g9754;
wire g3425;
wire II10135;
wire II7716;
wire g6397;
wire II13203;
wire g6689;
wire II8418;
wire II5867;
wire g7775;
wire g11581;
wire g4377;
wire g8094;
wire g8076;
wire II16920;
wire g11510;
wire g10555;
wire g6178;
wire II5295;
wire g8389;
wire II12904;
wire g4193;
wire g5212;
wire g9887;
wire g10589;
wire g5690;
wire II5613;
wire g7309;
wire II13197;
wire II14961;
wire II14779;
wire II7240;
wire g3537;
wire II9875;
wire g10368;
wire II13266;
wire II5025;
wire g7737;
wire g5034;
wire g2339;
wire II5672;
wire g10283;
wire g4498;
wire g7637;
wire g11348;
wire g3996;
wire g3519;
wire II9023;
wire g7706;
wire g2652;
wire g11384;
wire g11042;
wire g2069;
wire g7730;
wire g10500;
wire g11175;
wire g4879;
wire g6154;
wire g8615;
wire g4794;
wire II10144;
wire g2255;
wire II7559;
wire g6081;
wire II15807;
wire g7046;
wire g4191;
wire g11555;
wire g10161;
wire II17331;
wire II9365;
wire II15565;
wire II9539;
wire II8535;
wire II5342;
wire g5866;
wire II13877;
wire II13051;
wire II13436;
wire II17108;
wire g7473;
wire II15057;
wire g8674;
wire g8701;
wire g10156;
wire g2216;
wire g6348;
wire g6203;
wire II10659;
wire II17616;
wire g6482;
wire g5598;
wire g9746;
wire g98;
wire g8177;
wire g8748;
wire II7639;
wire g8656;
wire II14252;
wire g5591;
wire g10354;
wire g5700;
wire II15994;
wire g11084;
wire II8282;
wire g4262;
wire g8754;
wire g3098;
wire II16601;
wire II15082;
wire g6442;
wire II14112;
wire II5922;
wire II12436;
wire g8420;
wire g9653;
wire g5830;
wire g10643;
wire g7466;
wire g2007;
wire II8662;
wire g5081;
wire II10963;
wire II5591;
wire g6880;
wire g6463;
wire g5032;
wire g11085;
wire g2807;
wire II16956;
wire g6088;
wire II17503;
wire g4504;
wire g8194;
wire g9939;
wire g5671;
wire g10065;
wire g8627;
wire II16160;
wire g7687;
wire g8963;
wire g10111;
wire g5481;
wire II10183;
wire g2861;
wire g3086;
wire g2021;
wire II9544;
wire g2028;
wire g8929;
wire g11076;
wire II6952;
wire g10458;
wire g7627;
wire II15332;
wire g10327;
wire g6073;
wire g10534;
wire g3337;
wire II11836;
wire g8922;
wire g7384;
wire II15716;
wire g3707;
wire g11423;
wire g6750;
wire g6647;
wire g10775;
wire g7183;
wire g5072;
wire g3877;
wire g10041;
wire g11408;
wire II7435;
wire g5169;
wire g6694;
wire g4286;
wire g2946;
wire g6576;
wire g5039;
wire g11112;
wire g7782;
wire g2629;
wire g7029;
wire g2205;
wire g7773;
wire g3814;
wire g9852;
wire g9943;
wire II16017;
wire g8291;
wire g1964;
wire g5887;
wire II16065;
wire g7335;
wire g9430;
wire g8569;
wire g11264;
wire g9697;
wire g4079;
wire II9276;
wire g7231;
wire g3521;
wire II12427;
wire g6039;
wire g11638;
wire II8611;
wire II4886;
wire g10529;
wire II14973;
wire g10612;
wire g4440;
wire g8330;
wire g9418;
wire g10798;
wire g4872;
wire g6801;
wire g5285;
wire II4986;
wire g11098;
wire g9802;
wire g3752;
wire g2914;
wire g3528;
wire g5817;
wire g10856;
wire II9016;
wire g4971;
wire g5532;
wire g9365;
wire II16236;
wire g8339;
wire II10231;
wire g4771;
wire g4801;
wire II5248;
wire II7803;
wire II11915;
wire g6251;
wire g9270;
wire g3941;
wire II5430;
wire II6037;
wire g5225;
wire g3113;
wire II6815;
wire g5796;
wire II8750;
wire g2530;
wire g2731;
wire II7478;
wire g2259;
wire g6732;
wire g7954;
wire II6022;
wire g8818;
wire II12106;
wire II5283;
wire g3943;
wire g3736;
wire g6843;
wire g8358;
wire II14216;
wire g3688;
wire II14684;
wire g8203;
wire II6186;
wire g11610;
wire g10277;
wire g4082;
wire g2347;
wire II11937;
wire g9173;
wire g7541;
wire g9721;
wire II14903;
wire g7548;
wire g4765;
wire g5508;
wire g4425;
wire II4942;
wire II14203;
wire II15545;
wire g9340;
wire II15263;
wire g3698;
wire II15968;
wire II15878;
wire g3247;
wire g5826;
wire g9844;
wire g3582;
wire g8858;
wire II16859;
wire g11179;
wire g9819;
wire g2168;
wire II10643;
wire II16553;
wire g8484;
wire II6968;
wire g6323;
wire II15253;
wire II14424;
wire g10431;
wire g2745;
wire g8935;
wire II7280;
wire II17146;
wire g4530;
wire g7824;
wire g3635;
wire g10541;
wire II17387;
wire g9974;
wire II5710;
wire g6134;
wire II13531;
wire II7061;
wire g10168;
wire g11292;
wire g5249;
wire II14040;
wire g7561;
wire g10426;
wire g2643;
wire g9689;
wire g4913;
wire g4593;
wire g5479;
wire g5732;
wire g8429;
wire g4351;
wire g4520;
wire g5402;
wire g4256;
wire g4163;
wire g7302;
wire g7007;
wire g8512;
wire g8519;
wire g4935;
wire II11207;
wire g2772;
wire g6275;
wire g11412;
wire II9102;
wire g11505;
wire g11592;
wire II8827;
wire II13248;
wire g2617;
wire g4315;
wire g9816;
wire g3744;
wire II5357;
wire II6310;
wire g7242;
wire g10088;
wire g2363;
wire II16427;
wire g8387;
wire g6106;
wire g4734;
wire g5842;
wire g6326;
wire g5663;
wire g2047;
wire g8128;
wire g8002;
wire g3038;
wire g10875;
wire II11908;
wire g4251;
wire g7260;
wire II9147;
wire II9194;
wire II5892;
wire II6767;
wire g6272;
wire II12114;
wire g10736;
wire g8264;
wire g4780;
wire II5005;
wire g4727;
wire II15736;
wire g3977;
wire g4487;
wire II17246;
wire II11665;
wire II14415;
wire g8015;
wire II6040;
wire g6727;
wire g10691;
wire II5865;
wire II15443;
wire II15607;
wire g9840;
wire g8433;
wire g2325;
wire g4275;
wire g7063;
wire II13969;
wire II4928;
wire II10549;
wire g10898;
wire g10973;
wire g8283;
wire g8949;
wire II15775;
wire g7437;
wire II13415;
wire g11321;
wire II11155;
wire g5415;
wire II6007;
wire g10706;
wire II16032;
wire II6821;
wire g6433;
wire g5271;
wire g6559;
wire g9724;
wire g10885;
wire g3102;
wire g9641;
wire g10208;
wire II16416;
wire II7308;
wire g5115;
wire g7800;
wire g5771;
wire II7384;
wire g11308;
wire g7496;
wire II16467;
wire g2097;
wire II9658;
wire g8483;
wire II9588;
wire g4159;
wire g3747;
wire g6266;
wire II10186;
wire g8183;
wire II13529;
wire II5202;
wire g10242;
wire g11211;
wire II12245;
wire II5606;
wire g3544;
wire g8589;
wire II5126;
wire g10633;
wire g8450;
wire II9132;
wire g10098;
wire g3880;
wire II15554;
wire g10491;
wire g10314;
wire g4400;
wire II11119;
wire II13364;
wire g4921;
wire II12999;
wire g2635;
wire g4475;
wire II7390;
wire II10081;
wire g7764;
wire II12235;
wire g2276;
wire II15615;
wire g5586;
wire g2170;
wire g7807;
wire g5918;
wire g9812;
wire g4230;
wire g11027;
wire g8513;
wire g2895;
wire g2195;
wire g11542;
wire II15290;
wire II5098;
wire II15232;
wire g3722;
wire g8693;
wire g10744;
wire g9313;
wire g7444;
wire II10729;
wire II16439;
wire II7264;
wire g4894;
wire g8551;
wire II5549;
wire II6904;
wire g7240;
wire II11169;
wire g4060;
wire g9308;
wire g10664;
wire g11280;
wire g5291;
wire g7958;
wire g11153;
wire g5810;
wire g11151;
wire II9948;
wire g9865;
wire g3791;
wire g5278;
wire g9662;
wire g1972;
wire g7585;
wire g8298;
wire g11104;
wire g9994;
wire g5002;
wire g3214;
wire II8716;
wire g3563;
wire g9735;
wire II5332;
wire g6121;
wire II11638;
wire g10235;
wire g7501;
wire g6823;
wire II5035;
wire g9614;
wire II13895;
wire g8880;
wire II8275;
wire II13767;
wire g4122;
wire g10671;
wire g9587;
wire II8943;
wire II17395;
wire g5146;
wire II9427;
wire g7286;
wire g6545;
wire II7194;
wire II9886;
wire g6903;
wire II5198;
wire g2235;
wire g2919;
wire II8589;
wire II8967;
wire g11236;
wire g7630;
wire g7876;
wire g11602;
wire g4962;
wire II13726;
wire II16044;
wire g5876;
wire g10434;
wire g2011;
wire g7872;
wire g6740;
wire II13086;
wire g9516;
wire g9026;
wire II15801;
wire g5614;
wire II13505;
wire II8385;
wire g3307;
wire g2868;
wire g9968;
wire g6338;
wire g11479;
wire g6714;
wire g11444;
wire g5611;
wire g9918;
wire II5484;
wire II11578;
wire g7294;
wire g2310;
wire g5893;
wire II16843;
wire g4870;
wire II7076;
wire II16623;
wire g7649;
wire g2570;
wire g6759;
wire g6297;
wire II8669;
wire g8707;
wire g4672;
wire g8879;
wire II15177;
wire g4828;
wire II17377;
wire g8101;
wire II17736;
wire II15752;
wire II12162;
wire II14442;
wire g2249;
wire II15823;
wire g9912;
wire g8813;
wire II5494;
wire g8266;
wire II6088;
wire II12616;
wire g11036;
wire g6413;
wire II12799;
wire II15063;
wire II10495;
wire g5631;
wire g11578;
wire II6121;
wire II16023;
wire II4955;
wire II8647;
wire II13949;
wire g8148;
wire II14090;
wire g10563;
wire g2537;
wire II12255;
wire II10036;
wire II15977;
wire g6723;
wire II11082;
wire II5716;
wire II11982;
wire II13800;
wire g10514;
wire g9898;
wire II7536;
wire g2640;
wire II11198;
wire g8744;
wire II13448;
wire II8761;
wire g6257;
wire g6921;
wire g10142;
wire g8840;
wire g4563;
wire g4252;
wire II11932;
wire g7967;
wire g10421;
wire g6806;
wire g4483;
wire II12038;
wire g11571;
wire II8262;
wire g10477;
wire g3501;
wire II8880;
wire g9618;
wire II12690;
wire II5641;
wire II17698;
wire g9710;
wire g9779;
wire II12825;
wire g10149;
wire g7611;
wire g8181;
wire g4591;
wire g4534;
wire g4519;
wire II11950;
wire g7579;
wire g2795;
wire g9890;
wire g5803;
wire g11156;
wire g8599;
wire g7422;
wire g10127;
wire II9880;
wire II5887;
wire II5106;
wire g10293;
wire g4087;
wire g3344;
wire g8312;
wire g4200;
wire g11607;
wire II16717;
wire II4879;
wire g2817;
wire II14388;
wire II5470;
wire g8822;
wire g11394;
wire II6888;
wire II15551;
wire g8308;
wire g4130;
wire II6094;
wire g9719;
wire g6508;
wire g2424;
wire g2654;
wire g9600;
wire g8321;
wire g5652;
wire g4271;
wire g6317;
wire g7749;
wire g4806;
wire g5657;
wire g6907;
wire g9388;
wire g6163;
wire II13568;
wire II11575;
wire II8624;
wire g3397;
wire II10343;
wire g2904;
wire g8609;
wire g11354;
wire II15432;
wire g11432;
wire g2352;
wire g7845;
wire g4974;
wire g4768;
wire II12156;
wire II5600;
wire g10826;
wire g8244;
wire g7921;
wire II13609;
wire g5426;
wire g2905;
wire g7032;
wire g10551;
wire g5769;
wire g8146;
wire II17444;
wire II13975;
wire g6666;
wire g2514;
wire g4319;
wire II5976;
wire g2071;
wire g3096;
wire II7272;
wire g4452;
wire g6734;
wire g3304;
wire II10147;
wire II14642;
wire g5214;
wire g6737;
wire g2231;
wire g7311;
wire g6820;
wire g4375;
wire g8572;
wire g1963;
wire g5204;
wire II13580;
wire g7085;
wire g8042;
wire II9326;
wire g8472;
wire g4297;
wire II10045;
wire II6049;
wire g9362;
wire g10220;
wire II17381;
wire g6551;
wire g5572;
wire II13991;
wire g5042;
wire g2874;
wire II6898;
wire g7923;
wire II13048;
wire g4761;
wire II5304;
wire g9094;
wire g4990;
wire II5655;
wire g7994;
wire II9981;
wire g7035;
wire g9921;
wire II17209;
wire g2187;
wire II13382;
wire II7743;
wire g8179;
wire II15500;
wire g11054;
wire II12248;
wire g10719;
wire II9585;
wire II8854;
wire g11547;
wire g11024;
wire g7058;
wire II14570;
wire g5904;
wire II15368;
wire g7689;
wire II13908;
wire II14549;
wire g5522;
wire g4190;
wire II12936;
wire g5897;
wire II17290;
wire g11066;
wire g8346;
wire g6244;
wire II9491;
wire g7279;
wire II5218;
wire g8799;
wire II6145;
wire g10436;
wire g7323;
wire g7318;
wire II16577;
wire g6453;
wire g8847;
wire g5781;
wire II11656;
wire II17327;
wire II14418;
wire g11482;
wire II17173;
wire II12360;
wire gbuf14;
wire II7671;
wire II17710;
wire g10083;
wire g6786;
wire g7980;
wire g8993;
wire g9745;
wire g4776;
wire g2435;
wire g7819;
wire II11191;
wire g9412;
wire g7124;
wire g6928;
wire II16074;
wire II7140;
wire g8632;
wire II11560;
wire II17359;
wire g11166;
wire II11641;
wire g11458;
wire II13630;
wire II6611;
wire g7704;
wire II15792;
wire g8715;
wire g8286;
wire g11398;
wire g5190;
wire g3731;
wire II14799;
wire II6876;
wire g2501;
wire II10509;
wire g10486;
wire g8259;
wire g6835;
wire g7789;
wire II15305;
wire II8503;
wire g2871;
wire g9350;
wire g8292;
wire g9609;
wire g6717;
wire g9428;
wire g11460;
wire g3121;
wire g4102;
wire II13002;
wire g10074;
wire g6047;
wire II5592;
wire II15892;
wire II15899;
wire g8080;
wire II4850;
wire II8919;
wire g5646;
wire g3987;
wire g9855;
wire g9082;
wire g11011;
wire g2764;
wire II16528;
wire II11456;
wire II5128;
wire g4676;
wire g8078;
wire g4369;
wire g5124;
wire g10819;
wire II7468;
wire g8887;
wire II8298;
wire g5901;
wire g2528;
wire II12857;
wire II6565;
wire g7888;
wire II8729;
wire g3427;
wire g8353;
wire g8217;
wire II13956;
wire g6944;
wire II14364;
wire g6290;
wire g9769;
wire II4903;
wire g3765;
wire g8073;
wire g8973;
wire g3070;
wire g4523;
wire g10883;
wire g11226;
wire g10344;
wire g5556;
wire II8004;
wire II8779;
wire II13574;
wire g11187;
wire g4384;
wire g8992;
wire g10196;
wire II16793;
wire II15406;
wire II9332;
wire g7623;
wire II6370;
wire g11312;
wire g4320;
wire II6294;
wire g10171;
wire g7893;
wire g11427;
wire g7979;
wire g6585;
wire g5175;
wire g4902;
wire g9937;
wire g3009;
wire II5116;
wire g11497;
wire g7057;
wire g6098;
wire g2840;
wire g10781;
wire II16148;
wire g9666;
wire g4281;
wire II6461;
wire g4360;
wire g5685;
wire II10299;
wire II15733;
wire g6538;
wire II8528;
wire g4055;
wire II14101;
wire II15272;
wire II9759;
wire g10132;
wire g4754;
wire II11354;
wire g5557;
wire g3088;
wire II10991;
wire g3818;
wire II11255;
wire g8230;
wire g10358;
wire II16583;
wire II10917;
wire g8221;
wire g10476;
wire g9880;
wire g6027;
wire g10444;
wire g9655;
wire g7945;
wire II13538;
wire g10804;
wire g2942;
wire g3524;
wire g2949;
wire g6526;
wire g10909;
wire g2838;
wire g6548;
wire g6042;
wire g4554;
wire g9759;
wire II5804;
wire g9530;
wire g11376;
wire g10371;
wire II14607;
wire g6218;
wire g6916;
wire g4729;
wire II11309;
wire g6234;
wire g8440;
wire II9789;
wire II8479;
wire g5013;
wire II6109;
wire g8683;
wire g4544;
wire g4416;
wire g6791;
wire g4576;
wire II11752;
wire II16664;
wire g10623;
wire g9730;
wire g6180;
wire g7739;
wire II9766;
wire g5692;
wire g4968;
wire g9268;
wire g11449;
wire II5184;
wire g8554;
wire g3292;
wire II11140;
wire g7378;
wire g8545;
wire g2521;
wire g8098;
wire g4390;
wire g2309;
wire g11243;
wire g5543;
wire II12805;
wire g7343;
wire g6478;
wire g7934;
wire II15421;
wire II12843;
wire g5255;
wire g8734;
wire II15341;
wire g11301;
wire g5755;
wire II13308;
wire II13809;
wire g11147;
wire II17716;
wire g7917;
wire g10118;
wire II10840;
wire g11275;
wire g2109;
wire g5266;
wire II7916;
wire g6399;
wire II10114;
wire II14582;
wire II5754;
wire II6432;
wire g11252;
wire II11472;
wire II14944;
wire II9475;
wire g5229;
wire II11605;
wire II10663;
wire II7586;
wire II17424;
wire II4869;
wire g6564;
wire g6403;
wire g4942;
wire g3461;
wire II13741;
wire g5007;
wire g6860;
wire II15350;
wire II15371;
wire g8773;
wire g7369;
wire II13825;
wire g5023;
wire g10178;
wire g2102;
wire II5229;
wire g5272;
wire g2478;
wire II14188;
wire g11465;
wire g8326;
wire g4098;
wire g5144;
wire g6002;
wire g4615;
wire g7088;
wire g2937;
wire g6627;
wire II7685;
wire II9359;
wire II6760;
wire II12271;
wire II17534;
wire g5195;
wire g3061;
wire II6844;
wire II14503;
wire g9505;
wire g3348;
wire II11716;
wire II9074;
wire g5063;
wire g6887;
wire II12942;
wire g8405;
wire g7415;
wire g5998;
wire II8442;
wire g8950;
wire II13907;
wire g2380;
wire g7970;
wire g10595;
wire II8421;
wire g10388;
wire g7740;
wire g6948;
wire g5728;
wire g5320;
wire g6285;
wire g6638;
wire g6811;
wire II10937;
wire II13418;
wire II12553;
wire g7116;
wire II16292;
wire g4836;
wire g11451;
wire g2348;
wire g8770;
wire II11997;
wire II17613;
wire g6192;
wire g6195;
wire II10825;
wire II14409;
wire g2080;
wire g4586;
wire II9744;
wire g3714;
wire g7910;
wire g5348;
wire II17666;
wire g3411;
wire g11317;
wire II13427;
wire g8726;
wire g6501;
wire g8093;
wire II7782;
wire II11498;
wire g8300;
wire II5230;
wire g10184;
wire II9594;
wire g3439;
wire g3418;
wire g5493;
wire g5699;
wire g4344;
wire g7077;
wire II5949;
wire g2224;
wire II13466;
wire g11341;
wire g2341;
wire g4330;
wire II12335;
wire g7580;
wire g9878;
wire II5406;
wire g10313;
wire g9949;
wire II6929;
wire II17116;
wire g11283;
wire II17315;
wire g5534;
wire g8337;
wire II14319;
wire g9423;
wire g11417;
wire g8270;
wire g7333;
wire g10509;
wire g3546;
wire g11294;
wire g7674;
wire g8792;
wire g10767;
wire g6161;
wire g10266;
wire g2912;
wire II17707;
wire g10796;
wire II4992;
wire g6061;
wire II17274;
wire g4773;
wire g10249;
wire II10314;
wire g4976;
wire g9923;
wire g9510;
wire g5885;
wire II16030;
wire g10848;
wire II16206;
wire g11636;
wire II6484;
wire II13023;
wire II16009;
wire II16673;
wire g6037;
wire g4077;
wire g7300;
wire g10257;
wire II13893;
wire II14218;
wire g6852;
wire g8028;
wire g5113;
wire II6071;
wire g4462;
wire g3738;
wire II10362;
wire II10427;
wire g11106;
wire II5060;
wire II13274;
wire g5097;
wire g3637;
wire g9699;
wire II13424;
wire g6578;
wire g3908;
wire II9706;
wire g8153;
wire g6918;
wire II15494;
wire g4442;
wire II11483;
wire g4084;
wire g3749;
wire g8411;
wire II4965;
wire g2159;
wire g2449;
wire II17362;
wire II15741;
wire g5625;
wire II13782;
wire II8050;
wire II17219;
wire II17767;
wire g8199;
wire g9024;
wire II15068;
wire II10296;
wire g3430;
wire g6935;
wire g8538;
wire g6633;
wire g8805;
wire g7133;
wire g11648;
wire g2888;
wire II14567;
wire II12493;
wire II12448;
wire g7478;
wire g11064;
wire g2247;
wire g11177;
wire g5083;
wire II14323;
wire g2317;
wire II13606;
wire g6889;
wire II13819;
wire II11391;
wire II14191;
wire g9324;
wire II11680;
wire g10567;
wire II16778;
wire g2250;
wire II7202;
wire g10116;
wire II16850;
wire II6150;
wire II14477;
wire g7515;
wire g4392;
wire g8567;
wire II15562;
wire II10762;
wire g10093;
wire II16025;
wire g5911;
wire II8641;
wire II8061;
wire g4089;
wire g9885;
wire II12523;
wire g7912;
wire II16283;
wire g10590;
wire g11303;
wire II11046;
wire g4473;
wire g5404;
wire g9535;
wire II5186;
wire II12208;
wire g3879;
wire g2040;
wire II7694;
wire g2191;
wire II15210;
wire II14939;
wire II15114;
wire II15993;
wire II16685;
wire g5036;
wire g8751;
wire g5647;
wire g8285;
wire g6891;
wire II10378;
wire II7043;
wire g10163;
wire g5501;
wire g3372;
wire g6808;
wire II10837;
wire g2481;
wire II13057;
wire g5844;
wire II8770;
wire g4268;
wire g11173;
wire II9114;
wire g4747;
wire g2218;
wire g6856;
wire II10204;
wire g8085;
wire II5137;
wire g6246;
wire g3254;
wire g5472;
wire g7072;
wire g8007;
wire II12565;
wire g10381;
wire g8351;
wire g4890;
wire g11044;
wire g9454;
wire g4581;
wire g3566;
wire g6418;
wire II12322;
wire g10891;
wire g6096;
wire g6831;
wire g2863;
wire g10198;
wire g4317;
wire II9084;
wire II14358;
wire g11082;
wire g8422;
wire II12040;
wire g11429;
wire II8179;
wire II12202;
wire g11553;
wire II12631;
wire g8988;
wire g7735;
wire II15299;
wire g6595;
wire II10613;
wire II17456;
wire g10336;
wire II12418;
wire II9296;
wire II13633;
wire g5483;
wire g5167;
wire g4787;
wire g2991;
wire g4602;
wire g10773;
wire g7027;
wire g10532;
wire II17540;
wire g3974;
wire II6289;
wire II7810;
wire g5361;
wire II9608;
wire II7746;
wire g7952;
wire II10910;
wire II6694;
wire g9826;
wire g9204;
wire II17092;
wire II13887;
wire g2200;
wire g7435;
wire g11420;
wire g9770;
wire g2257;
wire g7793;
wire g2169;
wire II5461;
wire g6649;
wire g10445;
wire g6209;
wire g5898;
wire g10285;
wire g8279;
wire II16124;
wire II6601;
wire g6304;
wire II13788;
wire g10859;
wire II4979;
wire g3050;
wire II11734;
wire g7811;
wire II10006;
wire g11323;
wire g8192;
wire II17390;
wire g6653;
wire g7919;
wire II8515;
wire g2337;
wire g9110;
wire g7464;
wire g9266;
wire g2023;
wire g5539;
wire g4234;
wire II11079;
wire g7471;
wire II13451;
wire g7762;
wire g10931;
wire g4288;
wire g5640;
wire g3709;
wire II12421;
wire g10057;
wire II5517;
wire g8942;
wire g4469;
wire g6292;
wire g11074;
wire g11091;
wire g5891;
wire g7771;
wire II9268;
wire g5588;
wire g4358;
wire g4496;
wire g8927;
wire g9592;
wire g3108;
wire g9589;
wire II15718;
wire g5809;
wire g9668;
wire g7525;
wire g6873;
wire g5783;
wire II11363;
wire g7559;
wire II15829;
wire g2707;
wire g7272;
wire II10078;
wire g8650;
wire g7503;
wire g4892;
wire II4911;
wire g7620;
wire g8465;
wire g6146;
wire g6772;
wire g10946;
wire II10289;
wire g2154;
wire g8811;
wire II16432;
wire g11549;
wire g4869;
wire g3694;
wire g7446;
wire II7166;
wire g7550;
wire g4165;
wire II11103;
wire g10211;
wire g9359;
wire II9346;
wire g9733;
wire II15238;
wire g9693;
wire II17746;
wire g5490;
wire II15675;
wire II10177;
wire II7022;
wire g6882;
wire g8548;
wire g10673;
wire II12433;
wire g3305;
wire g7659;
wire g3798;
wire II6316;
wire II15224;
wire g5616;
wire g10237;
wire g7843;
wire g4242;
wire g9356;
wire II10105;
wire g2725;
wire g1974;
wire g6030;
wire g9416;
wire g7852;
wire g3388;
wire II14701;
wire g4260;
wire g11653;
wire g5000;
wire g8624;
wire II9988;
wire g9291;
wire II10949;
wire g8136;
wire g4822;
wire II7322;
wire II6587;
wire g4867;
wire g9085;
wire g10120;
wire g8268;
wire g8838;
wire g4908;
wire g8103;
wire g8933;
wire II12067;
wire II16039;
wire II6200;
wire II11707;
wire g10139;
wire II6302;
wire g5354;
wire g6833;
wire II5540;
wire g8705;
wire II16356;
wire g2809;
wire g6349;
wire g8746;
wire g8731;
wire g5301;
wire g7798;
wire II15665;
wire g5596;
wire g11228;
wire g4529;
wire II9421;
wire g3727;
wire II17237;
wire g6411;
wire g8696;
wire g10539;
wire II7546;
wire g2540;
wire g2077;
wire g9954;
wire g3012;
wire g3624;
wire II8465;
wire g2851;
wire II8872;
wire g6539;
wire g9780;
wire g11164;
wire II7952;
wire g2508;
wire g3910;
wire g9346;
wire g7292;
wire g4224;
wire g7572;
wire g6813;
wire II14232;
wire g4143;
wire g2304;
wire II8231;
wire g3793;
wire g6905;
wire g6671;
wire g3219;
wire g3800;
wire g2948;
wire II8109;
wire II5418;
wire g6344;
wire II14394;
wire g3101;
wire g8506;
wire g9910;
wire II9153;
wire g4223;
wire g10130;
wire g3998;
wire g11282;
wire II15317;
wire g5188;
wire g4886;
wire g4674;
wire g11576;
wire g4124;
wire II9108;
wire II13615;
wire II11746;
wire II10819;
wire g6331;
wire g3975;
wire g6104;
wire g10488;
wire II16525;
wire g10129;
wire II6746;
wire II11183;
wire II11901;
wire II12015;
wire g10683;
wire g4215;
wire II10248;
wire II5555;
wire g6328;
wire II5276;
wire g11495;
wire g6053;
wire g10788;
wire g7299;
wire g6043;
wire II15184;
wire g4278;
wire g5665;
wire g4431;
wire g7693;
wire g10322;
wire II10855;
wire II5879;
wire g11560;
wire g9814;
wire II15442;
wire g8956;
wire g5181;
wire II15437;
wire g3204;
wire g5317;
wire II5880;
wire g10933;
wire II10171;
wire g8262;
wire g2162;
wire g6354;
wire g7542;
wire II7182;
wire g6072;
wire II14602;
wire II15832;
wire II5475;
wire g6016;
wire g9952;
wire II7029;
wire g6532;
wire g7618;
wire g2829;
wire g10734;
wire II12981;
wire g6757;
wire g4049;
wire g4782;
wire g2297;
wire g4171;
wire g4273;
wire II9712;
wire g11641;
wire g2951;
wire II11662;
wire g5707;
wire g7597;
wire g8126;
wire g4166;
wire II12035;
wire g5938;
wire II8473;
wire II11569;
wire g7257;
wire g5088;
wire g9604;
wire g6270;
wire g7414;
wire g5103;
wire g4485;
wire II5435;
wire II15971;
wire g4438;
wire g10873;
wire g8408;
wire g9648;
wire g5296;
wire g7122;
wire g4875;
wire II5704;
wire II11692;
wire g9942;
wire II15204;
wire II14614;
wire g3111;
wire g9984;
wire II5324;
wire g8870;
wire g2031;
wire g6388;
wire g8920;
wire g9657;
wire II14299;
wire II15430;
wire g3227;
wire g6581;
wire II5571;
wire g5702;
wire II6133;
wire g4557;
wire g6719;
wire g3381;
wire g7245;
wire g6749;
wire II6679;
wire II9138;
wire g6079;
wire II16053;
wire g4381;
wire g7533;
wire II13284;
wire g2620;
wire II5824;
wire g8515;
wire II10810;
wire II9995;
wire g6845;
wire II17585;
wire II14713;
wire g4112;
wire g8481;
wire g11198;
wire II5695;
wire g6119;
wire II15701;
wire g10701;
wire g3979;
wire II7054;
wire II17555;
wire II7224;
wire II13485;
wire g9620;
wire g8498;
wire g11025;
wire g2638;
wire g2197;
wire g7759;
wire g2756;
wire g4680;
wire g4450;
wire II15075;
wire g10240;
wire II16037;
wire II9180;
wire II9773;
wire g5942;
wire g8947;
wire II5445;
wire II13965;
wire g2779;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g30 <= 0;
  else
    g30 <= g6254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g31 <= 0;
  else
    g31 <= g6255;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g32 <= 0;
  else
    g32 <= g11397;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g33 <= 0;
  else
    g33 <= g10867;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g34 <= 0;
  else
    g34 <= g10868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g35 <= 0;
  else
    g35 <= g10869;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g36 <= 0;
  else
    g36 <= g10870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g37 <= 0;
  else
    g37 <= g10871;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g38 <= 0;
  else
    g38 <= g10872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g39 <= 0;
  else
    g39 <= g10774;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g40 <= 0;
  else
    g40 <= g10775;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g41 <= 0;
  else
    g41 <= g6256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g42 <= 0;
  else
    g42 <= g6257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g43 <= 0;
  else
    g43 <= g6258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g44 <= 0;
  else
    g44 <= g6259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g45 <= 0;
  else
    g45 <= g6260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g46 <= 0;
  else
    g46 <= g6261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g47 <= 0;
  else
    g47 <= g6262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g48 <= 0;
  else
    g48 <= g6263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g82 <= 0;
  else
    g82 <= g6264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g83 <= 0;
  else
    g83 <= g6265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g84 <= 0;
  else
    g84 <= g6266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g85 <= 0;
  else
    g85 <= g6267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g86 <= 0;
  else
    g86 <= g6268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g87 <= 0;
  else
    g87 <= g6269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g88 <= 0;
  else
    g88 <= g6270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g89 <= 0;
  else
    g89 <= g6271;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g90 <= 0;
  else
    g90 <= g6272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g91 <= 0;
  else
    g91 <= g6273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g92 <= 0;
  else
    g92 <= g6274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g93 <= 0;
  else
    g93 <= g6275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g94 <= 0;
  else
    g94 <= g6276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g95 <= 0;
  else
    g95 <= g6277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g96 <= 0;
  else
    g96 <= g6278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g99 <= 0;
  else
    g99 <= g6279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g100 <= 0;
  else
    g100 <= g6280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g101 <= 0;
  else
    g101 <= g6281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g102 <= 0;
  else
    g102 <= g6282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g103 <= 0;
  else
    g103 <= g6283;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g104 <= 0;
  else
    g104 <= g6284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g28 <= 0;
  else
    g28 <= g6285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g29 <= 0;
  else
    g29 <= g6253;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g898 <= 0;
  else
    g898 <= g4195;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g901 <= 0;
  else
    g901 <= g4197;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g904 <= 0;
  else
    g904 <= g4198;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g907 <= 0;
  else
    g907 <= g4199;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g910 <= 0;
  else
    g910 <= g4200;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g913 <= 0;
  else
    g913 <= g4201;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g916 <= 0;
  else
    g916 <= g4202;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g919 <= 0;
  else
    g919 <= g4203;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g922 <= 0;
  else
    g922 <= g4204;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g925 <= 0;
  else
    g925 <= g4196;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g971 <= 0;
  else
    g971 <= g11470;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g976 <= 0;
  else
    g976 <= g11471;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g981 <= 0;
  else
    g981 <= g11472;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g986 <= 0;
  else
    g986 <= g11473;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g944 <= 0;
  else
    g944 <= g11398;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g947 <= 0;
  else
    g947 <= g11399;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g950 <= 0;
  else
    g950 <= g11400;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g953 <= 0;
  else
    g953 <= g11401;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g956 <= 0;
  else
    g956 <= g11402;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g959 <= 0;
  else
    g959 <= g11403;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g962 <= 0;
  else
    g962 <= g11404;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g965 <= 0;
  else
    g965 <= g11405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g968 <= 0;
  else
    g968 <= g11406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g886 <= 0;
  else
    g886 <= g4191;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g889 <= 0;
  else
    g889 <= g4192;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g892 <= 0;
  else
    g892 <= g4193;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g895 <= 0;
  else
    g895 <= g4194;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g928 <= 0;
  else
    g928 <= g8569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g932 <= 0;
  else
    g932 <= g8570;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g936 <= 0;
  else
    g936 <= g8571;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g940 <= 0;
  else
    g940 <= g8572;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g883 <= 0;
  else
    g883 <= g4897;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g882 <= 0;
  else
    g882 <= gbuf1;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g878 <= 0;
  else
    g878 <= g4896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g876 <= 0;
  else
    g876 <= gbuf2;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g757 <= 0;
  else
    g757 <= g11179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g755 <= 0;
  else
    g755 <= g6298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g756 <= 0;
  else
    g756 <= gbuf3;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g745 <= 0;
  else
    g745 <= g2639;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g746 <= 0;
  else
    g746 <= g2638;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g750 <= 0;
  else
    g750 <= g4171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g754 <= 0;
  else
    g754 <= g4895;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g758 <= 0;
  else
    g758 <= g6797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g762 <= 0;
  else
    g762 <= g6798;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g766 <= 0;
  else
    g766 <= g6799;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g770 <= 0;
  else
    g770 <= g7288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g774 <= 0;
  else
    g774 <= g7785;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g778 <= 0;
  else
    g778 <= g8076;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g782 <= 0;
  else
    g782 <= g8273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g786 <= 0;
  else
    g786 <= g8436;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g790 <= 0;
  else
    g790 <= g8567;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g865 <= 0;
  else
    g865 <= g8275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g794 <= 0;
  else
    g794 <= g6800;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g798 <= 0;
  else
    g798 <= g6801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g802 <= 0;
  else
    g802 <= g6802;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g806 <= 0;
  else
    g806 <= g7289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g810 <= 0;
  else
    g810 <= g7786;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g814 <= 0;
  else
    g814 <= g8077;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g818 <= 0;
  else
    g818 <= g8274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g822 <= 0;
  else
    g822 <= g8437;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g826 <= 0;
  else
    g826 <= g8568;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g829 <= 0;
  else
    g829 <= g4182;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g833 <= 0;
  else
    g833 <= g4183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g837 <= 0;
  else
    g837 <= g4184;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g841 <= 0;
  else
    g841 <= g4185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g845 <= 0;
  else
    g845 <= g4186;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g849 <= 0;
  else
    g849 <= g4187;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g853 <= 0;
  else
    g853 <= g4188;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g857 <= 0;
  else
    g857 <= g4189;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g861 <= 0;
  else
    g861 <= g4190;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g874 <= 0;
  else
    g874 <= g9821;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g868 <= 0;
  else
    g868 <= gbuf4;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g875 <= 0;
  else
    g875 <= g9822;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g869 <= 0;
  else
    g869 <= gbuf5;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g590 <= 0;
  else
    g590 <= g5653;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g584 <= 0;
  else
    g584 <= g6292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g585 <= 0;
  else
    g585 <= g6293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g586 <= 0;
  else
    g586 <= g6294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g587 <= 0;
  else
    g587 <= g6295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g588 <= 0;
  else
    g588 <= g6296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g589 <= 0;
  else
    g589 <= g6297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g578 <= 0;
  else
    g578 <= g6286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g579 <= 0;
  else
    g579 <= g6287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g580 <= 0;
  else
    g580 <= g6288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g581 <= 0;
  else
    g581 <= g6289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g582 <= 0;
  else
    g582 <= g6290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g583 <= 0;
  else
    g583 <= g6291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g253 <= 0;
  else
    g253 <= g7750;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g256 <= 0;
  else
    g256 <= g7752;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g257 <= 0;
  else
    g257 <= g7753;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g258 <= 0;
  else
    g258 <= g7754;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g259 <= 0;
  else
    g259 <= g7755;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g260 <= 0;
  else
    g260 <= g7756;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g261 <= 0;
  else
    g261 <= g7757;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g262 <= 0;
  else
    g262 <= g7758;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g254 <= 0;
  else
    g254 <= g7759;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g255 <= 0;
  else
    g255 <= g7751;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g143 <= 0;
  else
    g143 <= g7746;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g166 <= 0;
  else
    g166 <= g7747;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g139 <= 0;
  else
    g139 <= g8418;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g135 <= 0;
  else
    g135 <= g8419;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g131 <= 0;
  else
    g131 <= g8420;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g127 <= 0;
  else
    g127 <= g8421;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g170 <= 0;
  else
    g170 <= g8422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g174 <= 0;
  else
    g174 <= g8423;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g162 <= 0;
  else
    g162 <= g8424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g158 <= 0;
  else
    g158 <= g8425;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g153 <= 0;
  else
    g153 <= g8426;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g148 <= 0;
  else
    g148 <= g8427;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g178 <= 0;
  else
    g178 <= g7748;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g182 <= 0;
  else
    g182 <= g7749;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g126 <= 0;
  else
    g126 <= g5642;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g263 <= 0;
  else
    g263 <= g7760;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g266 <= 0;
  else
    g266 <= g7761;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g269 <= 0;
  else
    g269 <= g7762;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g272 <= 0;
  else
    g272 <= g7763;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g275 <= 0;
  else
    g275 <= g7764;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g278 <= 0;
  else
    g278 <= g7765;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g281 <= 0;
  else
    g281 <= g7766;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g284 <= 0;
  else
    g284 <= g7767;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g287 <= 0;
  else
    g287 <= g7768;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g290 <= 0;
  else
    g290 <= g7769;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g293 <= 0;
  else
    g293 <= g7770;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g296 <= 0;
  else
    g296 <= g7771;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g299 <= 0;
  else
    g299 <= g7772;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g302 <= 0;
  else
    g302 <= g7773;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g123 <= 0;
  else
    g123 <= g8272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g119 <= 0;
  else
    g119 <= g7745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g611 <= 0;
  else
    g611 <= g9930;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g617 <= 0;
  else
    g617 <= g8780;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g591 <= 0;
  else
    g591 <= g9818;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g599 <= 0;
  else
    g599 <= g9819;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g605 <= 0;
  else
    g605 <= g9820;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g630 <= 0;
  else
    g630 <= g7287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g631 <= 0;
  else
    g631 <= g5654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g632 <= 0;
  else
    g632 <= g5655;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g635 <= 0;
  else
    g635 <= g5656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g627 <= 0;
  else
    g627 <= g5657;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g636 <= 0;
  else
    g636 <= g8781;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g639 <= 0;
  else
    g639 <= g8063;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g622 <= 0;
  else
    g622 <= g9338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g643 <= 0;
  else
    g643 <= g8064;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g646 <= 0;
  else
    g646 <= g8065;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g650 <= 0;
  else
    g650 <= g8066;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g654 <= 0;
  else
    g654 <= g8067;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g658 <= 0;
  else
    g658 <= g9339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g668 <= 0;
  else
    g668 <= g9340;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g677 <= 0;
  else
    g677 <= g9341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g686 <= 0;
  else
    g686 <= g9342;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g695 <= 0;
  else
    g695 <= g9343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g704 <= 0;
  else
    g704 <= g9344;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g713 <= 0;
  else
    g713 <= g9345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g722 <= 0;
  else
    g722 <= g9346;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g731 <= 0;
  else
    g731 <= g9347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g664 <= 0;
  else
    g664 <= g8782;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g673 <= 0;
  else
    g673 <= g8428;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g682 <= 0;
  else
    g682 <= g8429;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g691 <= 0;
  else
    g691 <= g8430;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g700 <= 0;
  else
    g700 <= g8431;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g709 <= 0;
  else
    g709 <= g8432;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g718 <= 0;
  else
    g718 <= g8433;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g727 <= 0;
  else
    g727 <= g8434;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g736 <= 0;
  else
    g736 <= g8435;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g8 <= 0;
  else
    g8 <= g2613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g17 <= 0;
  else
    g17 <= g4894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g481 <= 0;
  else
    g481 <= g11324;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g486 <= 0;
  else
    g486 <= g11331;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g491 <= 0;
  else
    g491 <= g11332;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g496 <= 0;
  else
    g496 <= g11333;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g501 <= 0;
  else
    g501 <= g11334;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g506 <= 0;
  else
    g506 <= g11335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g511 <= 0;
  else
    g511 <= g11336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g516 <= 0;
  else
    g516 <= g11337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g476 <= 0;
  else
    g476 <= g11338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g542 <= 0;
  else
    g542 <= g11325;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g538 <= 0;
  else
    g538 <= g11326;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g534 <= 0;
  else
    g534 <= g11327;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g530 <= 0;
  else
    g530 <= g11328;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g525 <= 0;
  else
    g525 <= g11329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g521 <= 0;
  else
    g521 <= g11330;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g456 <= 0;
  else
    g456 <= g11466;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g461 <= 0;
  else
    g461 <= g11467;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g466 <= 0;
  else
    g466 <= g11468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g471 <= 0;
  else
    g471 <= g11469;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g305 <= 0;
  else
    g305 <= g5643;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g315 <= 0;
  else
    g315 <= g5645;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g318 <= 0;
  else
    g318 <= g5646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g321 <= 0;
  else
    g321 <= g5647;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g324 <= 0;
  else
    g324 <= g5648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g327 <= 0;
  else
    g327 <= g5649;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g330 <= 0;
  else
    g330 <= g5650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g333 <= 0;
  else
    g333 <= g5651;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g309 <= 0;
  else
    g309 <= g5652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g312 <= 0;
  else
    g312 <= g5644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g426 <= 0;
  else
    g426 <= g11256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g386 <= 0;
  else
    g386 <= g11263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g391 <= 0;
  else
    g391 <= g11264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g396 <= 0;
  else
    g396 <= g11265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g401 <= 0;
  else
    g401 <= g11266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g406 <= 0;
  else
    g406 <= g11267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g411 <= 0;
  else
    g411 <= g11268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g416 <= 0;
  else
    g416 <= g11269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g421 <= 0;
  else
    g421 <= g11270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g452 <= 0;
  else
    g452 <= g11257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g448 <= 0;
  else
    g448 <= g11258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g444 <= 0;
  else
    g444 <= g11259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g440 <= 0;
  else
    g440 <= g11260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g435 <= 0;
  else
    g435 <= g11261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g431 <= 0;
  else
    g431 <= g11262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g369 <= 0;
  else
    g369 <= g11439;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g374 <= 0;
  else
    g374 <= g11440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g378 <= 0;
  else
    g378 <= g11441;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g382 <= 0;
  else
    g382 <= g11442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g336 <= 0;
  else
    g336 <= g11653;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g348 <= 0;
  else
    g348 <= g11506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g351 <= 0;
  else
    g351 <= g11507;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g354 <= 0;
  else
    g354 <= g11508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g357 <= 0;
  else
    g357 <= g11509;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g360 <= 0;
  else
    g360 <= g11510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g363 <= 0;
  else
    g363 <= g11511;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g366 <= 0;
  else
    g366 <= g11512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g342 <= 0;
  else
    g342 <= g11513;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g339 <= 0;
  else
    g339 <= g11505;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g345 <= 0;
  else
    g345 <= g11642;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g49 <= 0;
  else
    g49 <= g7774;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g52 <= 0;
  else
    g52 <= g7777;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g55 <= 0;
  else
    g55 <= g7778;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g58 <= 0;
  else
    g58 <= g7779;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g61 <= 0;
  else
    g61 <= g7780;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g64 <= 0;
  else
    g64 <= g7781;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g67 <= 0;
  else
    g67 <= g7782;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g70 <= 0;
  else
    g70 <= g7783;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g73 <= 0;
  else
    g73 <= g7784;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g76 <= 0;
  else
    g76 <= g7775;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g79 <= 0;
  else
    g79 <= g7776;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g113 <= 0;
  else
    g113 <= g7285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g114 <= 0;
  else
    g114 <= gbuf6;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1955 <= 0;
  else
    g1955 <= g6338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1956 <= 0;
  else
    g1956 <= gbuf7;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1957 <= 0;
  else
    g1957 <= gbuf8;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1700 <= 0;
  else
    g1700 <= gbuf9;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1696 <= 0;
  else
    g1696 <= g6842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1703 <= 0;
  else
    g1703 <= g6843;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1710 <= 0;
  else
    g1710 <= g4901;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1713 <= 0;
  else
    g1713 <= g6336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1718 <= 0;
  else
    g1718 <= g6337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1766 <= 0;
  else
    g1766 <= g7810;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1771 <= 0;
  else
    g1771 <= g7811;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1776 <= 0;
  else
    g1776 <= g7812;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1781 <= 0;
  else
    g1781 <= g7813;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1786 <= 0;
  else
    g1786 <= g7814;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1791 <= 0;
  else
    g1791 <= g8080;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1796 <= 0;
  else
    g1796 <= g8280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1801 <= 0;
  else
    g1801 <= g8450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1806 <= 0;
  else
    g1806 <= g8573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1711 <= 0;
  else
    g1711 <= g6335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1834 <= 0;
  else
    g1834 <= g9895;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1840 <= 0;
  else
    g1840 <= g8694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1814 <= 0;
  else
    g1814 <= g9825;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1822 <= 0;
  else
    g1822 <= g9826;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1828 <= 0;
  else
    g1828 <= g9827;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1848 <= 0;
  else
    g1848 <= g7366;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1849 <= 0;
  else
    g1849 <= g5670;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1850 <= 0;
  else
    g1850 <= g5671;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1853 <= 0;
  else
    g1853 <= g5672;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1845 <= 0;
  else
    g1845 <= g5673;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1854 <= 0;
  else
    g1854 <= g11408;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1857 <= 0;
  else
    g1857 <= g11409;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1861 <= 0;
  else
    g1861 <= g7815;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1864 <= 0;
  else
    g1864 <= g7816;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1868 <= 0;
  else
    g1868 <= g7817;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1872 <= 0;
  else
    g1872 <= g9348;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1882 <= 0;
  else
    g1882 <= g9349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1891 <= 0;
  else
    g1891 <= g9350;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1900 <= 0;
  else
    g1900 <= g9351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1909 <= 0;
  else
    g1909 <= g9352;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1918 <= 0;
  else
    g1918 <= g9353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1927 <= 0;
  else
    g1927 <= g9354;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1936 <= 0;
  else
    g1936 <= g9355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1945 <= 0;
  else
    g1945 <= g9356;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1878 <= 0;
  else
    g1878 <= g8695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1887 <= 0;
  else
    g1887 <= g8281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1896 <= 0;
  else
    g1896 <= g8282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1905 <= 0;
  else
    g1905 <= g8283;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1914 <= 0;
  else
    g1914 <= g8284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1923 <= 0;
  else
    g1923 <= g8285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1932 <= 0;
  else
    g1932 <= g8286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1941 <= 0;
  else
    g1941 <= g8287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1950 <= 0;
  else
    g1950 <= g8288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g16 <= 0;
  else
    g16 <= g4906;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g7 <= 0;
  else
    g7 <= g2731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1736 <= 0;
  else
    g1736 <= g6846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1737 <= 0;
  else
    g1737 <= gbuf10;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1648 <= 0;
  else
    g1648 <= g11181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1651 <= 0;
  else
    g1651 <= g11182;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1642 <= 0;
  else
    g1642 <= g11183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1645 <= 0;
  else
    g1645 <= g11184;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1610 <= 0;
  else
    g1610 <= g6845;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1765 <= 0;
  else
    g1765 <= g3329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1811 <= 0;
  else
    g1811 <= g11185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1721 <= 0;
  else
    g1721 <= g10878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1724 <= 0;
  else
    g1724 <= g10879;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1727 <= 0;
  else
    g1727 <= g10880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1730 <= 0;
  else
    g1730 <= g10881;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1733 <= 0;
  else
    g1733 <= g10882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1738 <= 0;
  else
    g1738 <= g5661;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1741 <= 0;
  else
    g1741 <= g5662;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1744 <= 0;
  else
    g1744 <= g5663;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1747 <= 0;
  else
    g1747 <= g5664;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1750 <= 0;
  else
    g1750 <= g5665;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1753 <= 0;
  else
    g1753 <= g5666;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1756 <= 0;
  else
    g1756 <= g5667;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1759 <= 0;
  else
    g1759 <= g5668;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1762 <= 0;
  else
    g1762 <= g5669;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1958 <= 0;
  else
    g1958 <= g6339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1810 <= 0;
  else
    g1810 <= g2044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1959 <= 0;
  else
    g1959 <= g4217;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1707 <= 0;
  else
    g1707 <= g4907;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1690 <= 0;
  else
    g1690 <= g6844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1170 <= 0;
  else
    g1170 <= g4205;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1173 <= 0;
  else
    g1173 <= g4209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1176 <= 0;
  else
    g1176 <= g4210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1179 <= 0;
  else
    g1179 <= g4211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1182 <= 0;
  else
    g1182 <= g4212;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1185 <= 0;
  else
    g1185 <= g4213;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1188 <= 0;
  else
    g1188 <= g4214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1191 <= 0;
  else
    g1191 <= g4215;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1194 <= 0;
  else
    g1194 <= g4216;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1197 <= 0;
  else
    g1197 <= g4206;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1200 <= 0;
  else
    g1200 <= g4207;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1203 <= 0;
  else
    g1203 <= g4208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1169 <= 0;
  else
    g1169 <= g6314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g108 <= 0;
  else
    g108 <= g11593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1336 <= 0;
  else
    g1336 <= g11654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1341 <= 0;
  else
    g1341 <= g11655;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1346 <= 0;
  else
    g1346 <= g11656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1351 <= 0;
  else
    g1351 <= g11657;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1206 <= 0;
  else
    g1206 <= g4898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1361 <= 0;
  else
    g1361 <= gbuf11;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1360 <= 0;
  else
    g1360 <= g9824;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1216 <= 0;
  else
    g1216 <= gbuf12;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1217 <= 0;
  else
    g1217 <= g9823;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1212 <= 0;
  else
    g1212 <= gbuf13;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1209 <= 0;
  else
    g1209 <= g10873;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1215 <= 0;
  else
    g1215 <= g6315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1357 <= 0;
  else
    g1357 <= g6330;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1289 <= 0;
  else
    g1289 <= g5660;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1275 <= 0;
  else
    g1275 <= g11443;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1235 <= 0;
  else
    g1235 <= g7296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1240 <= 0;
  else
    g1240 <= g7297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1245 <= 0;
  else
    g1245 <= g7298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1250 <= 0;
  else
    g1250 <= g7299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1255 <= 0;
  else
    g1255 <= g7300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1260 <= 0;
  else
    g1260 <= g7301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1265 <= 0;
  else
    g1265 <= g7302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1270 <= 0;
  else
    g1270 <= g7303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1304 <= 0;
  else
    g1304 <= g7290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1300 <= 0;
  else
    g1300 <= g7291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1296 <= 0;
  else
    g1296 <= g7292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1292 <= 0;
  else
    g1292 <= g7293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1284 <= 0;
  else
    g1284 <= g7294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1280 <= 0;
  else
    g1280 <= g7295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1218 <= 0;
  else
    g1218 <= g8276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1223 <= 0;
  else
    g1223 <= g8277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1227 <= 0;
  else
    g1227 <= g8278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1231 <= 0;
  else
    g1231 <= g8279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1356 <= 0;
  else
    g1356 <= g6818;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1317 <= 0;
  else
    g1317 <= gbuf14;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1314 <= 0;
  else
    g1314 <= g11629;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1318 <= 0;
  else
    g1318 <= g11630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1321 <= 0;
  else
    g1321 <= g11631;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1324 <= 0;
  else
    g1324 <= g11632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1327 <= 0;
  else
    g1327 <= g11633;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1330 <= 0;
  else
    g1330 <= g11634;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1333 <= 0;
  else
    g1333 <= g11635;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1308 <= 0;
  else
    g1308 <= g11627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1311 <= 0;
  else
    g1311 <= g11628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1035 <= 0;
  else
    g1035 <= g7787;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1047 <= 0;
  else
    g1047 <= g7790;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1050 <= 0;
  else
    g1050 <= g7791;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1053 <= 0;
  else
    g1053 <= g7792;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1056 <= 0;
  else
    g1056 <= g7793;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1059 <= 0;
  else
    g1059 <= g7794;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1062 <= 0;
  else
    g1062 <= g7795;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1065 <= 0;
  else
    g1065 <= g7796;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1038 <= 0;
  else
    g1038 <= g7797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1041 <= 0;
  else
    g1041 <= g7788;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1044 <= 0;
  else
    g1044 <= g7789;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1068 <= 0;
  else
    g1068 <= g6803;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1080 <= 0;
  else
    g1080 <= g6806;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1083 <= 0;
  else
    g1083 <= g6807;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1086 <= 0;
  else
    g1086 <= g6808;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1089 <= 0;
  else
    g1089 <= g6809;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1092 <= 0;
  else
    g1092 <= g6810;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1095 <= 0;
  else
    g1095 <= g6811;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1098 <= 0;
  else
    g1098 <= g6812;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1074 <= 0;
  else
    g1074 <= g6813;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1071 <= 0;
  else
    g1071 <= g6804;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1077 <= 0;
  else
    g1077 <= g6805;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1027 <= 0;
  else
    g1027 <= g7798;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g995 <= 0;
  else
    g995 <= g7801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g991 <= 0;
  else
    g991 <= g7802;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1003 <= 0;
  else
    g1003 <= g7803;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g999 <= 0;
  else
    g999 <= g7804;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1011 <= 0;
  else
    g1011 <= g7805;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1007 <= 0;
  else
    g1007 <= g7806;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1019 <= 0;
  else
    g1019 <= g7807;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1015 <= 0;
  else
    g1015 <= g7808;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1023 <= 0;
  else
    g1023 <= g7799;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1032 <= 0;
  else
    g1032 <= g7800;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g105 <= 0;
  else
    g105 <= g11180;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1117 <= 0;
  else
    g1117 <= g6299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1121 <= 0;
  else
    g1121 <= g6306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1125 <= 0;
  else
    g1125 <= g6307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1129 <= 0;
  else
    g1129 <= g6308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1133 <= 0;
  else
    g1133 <= g6309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1137 <= 0;
  else
    g1137 <= g6310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1141 <= 0;
  else
    g1141 <= g6311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1145 <= 0;
  else
    g1145 <= g6312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1113 <= 0;
  else
    g1113 <= g6313;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1166 <= 0;
  else
    g1166 <= g6300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1163 <= 0;
  else
    g1163 <= g6301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1160 <= 0;
  else
    g1160 <= g6302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1157 <= 0;
  else
    g1157 <= g6303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1153 <= 0;
  else
    g1153 <= g6304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1149 <= 0;
  else
    g1149 <= g6305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1101 <= 0;
  else
    g1101 <= g6814;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1104 <= 0;
  else
    g1104 <= g6815;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1107 <= 0;
  else
    g1107 <= g6816;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1110 <= 0;
  else
    g1110 <= g6817;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1618 <= 0;
  else
    g1618 <= g11611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1615 <= 0;
  else
    g1615 <= g8868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1621 <= 0;
  else
    g1621 <= g8869;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1624 <= 0;
  else
    g1624 <= g8870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1627 <= 0;
  else
    g1627 <= g8871;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1630 <= 0;
  else
    g1630 <= g8872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1633 <= 0;
  else
    g1633 <= g8873;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1636 <= 0;
  else
    g1636 <= g8874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1639 <= 0;
  else
    g1639 <= g8448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1512 <= 0;
  else
    g1512 <= g8449;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1448 <= 0;
  else
    g1448 <= g11594;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1444 <= 0;
  else
    g1444 <= g8987;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1440 <= 0;
  else
    g1440 <= g8988;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1436 <= 0;
  else
    g1436 <= g8989;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1432 <= 0;
  else
    g1432 <= g8990;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1403 <= 0;
  else
    g1403 <= g8991;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1428 <= 0;
  else
    g1428 <= g8992;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1407 <= 0;
  else
    g1407 <= g8993;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1424 <= 0;
  else
    g1424 <= g7330;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1411 <= 0;
  else
    g1411 <= g7331;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1419 <= 0;
  else
    g1419 <= g7332;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1515 <= 0;
  else
    g1515 <= g7333;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1520 <= 0;
  else
    g1520 <= g7334;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1415 <= 0;
  else
    g1415 <= g7335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1453 <= 0;
  else
    g1453 <= g7326;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1458 <= 0;
  else
    g1458 <= g7327;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1462 <= 0;
  else
    g1462 <= g8438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1466 <= 0;
  else
    g1466 <= g8439;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1470 <= 0;
  else
    g1470 <= g8440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1474 <= 0;
  else
    g1474 <= g8441;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1478 <= 0;
  else
    g1478 <= g8442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1482 <= 0;
  else
    g1482 <= g8443;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1486 <= 0;
  else
    g1486 <= g8444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1490 <= 0;
  else
    g1490 <= g8445;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1494 <= 0;
  else
    g1494 <= g8446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1499 <= 0;
  else
    g1499 <= g8447;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1504 <= 0;
  else
    g1504 <= g7328;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1508 <= 0;
  else
    g1508 <= g7329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1393 <= 0;
  else
    g1393 <= g7320;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1394 <= 0;
  else
    g1394 <= g7809;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g115 <= 0;
  else
    g115 <= g7321;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g201 <= 0;
  else
    g201 <= g7304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1374 <= 0;
  else
    g1374 <= g6825;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g197 <= 0;
  else
    g197 <= g6835;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1389 <= 0;
  else
    g1389 <= g6836;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g192 <= 0;
  else
    g192 <= g6837;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1397 <= 0;
  else
    g1397 <= g7322;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g248 <= 0;
  else
    g248 <= g7323;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1400 <= 0;
  else
    g1400 <= g7324;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g243 <= 0;
  else
    g243 <= g7325;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1362 <= 0;
  else
    g1362 <= g7305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g237 <= 0;
  else
    g237 <= g7306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1365 <= 0;
  else
    g1365 <= g7307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g231 <= 0;
  else
    g231 <= g7319;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1368 <= 0;
  else
    g1368 <= g7308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g225 <= 0;
  else
    g225 <= g7309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1371 <= 0;
  else
    g1371 <= g7311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g219 <= 0;
  else
    g219 <= g7310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1377 <= 0;
  else
    g1377 <= g7312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g213 <= 0;
  else
    g213 <= g7313;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1380 <= 0;
  else
    g1380 <= g7314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g207 <= 0;
  else
    g207 <= g7315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1383 <= 0;
  else
    g1383 <= g7316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g186 <= 0;
  else
    g186 <= g7317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1386 <= 0;
  else
    g1386 <= g7318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4 <= 0;
  else
    g4 <= g8079;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g12 <= 0;
  else
    g12 <= g7337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1 <= 0;
  else
    g1 <= g8078;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g9 <= 0;
  else
    g9 <= g7336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1527 <= 0;
  else
    g1527 <= g4899;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1524 <= 0;
  else
    g1524 <= g7338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1528 <= 0;
  else
    g1528 <= g7339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1531 <= 0;
  else
    g1531 <= g7340;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1534 <= 0;
  else
    g1534 <= g7341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1537 <= 0;
  else
    g1537 <= g7342;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1540 <= 0;
  else
    g1540 <= g7343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1543 <= 0;
  else
    g1543 <= g7344;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1546 <= 0;
  else
    g1546 <= g7345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1549 <= 0;
  else
    g1549 <= g7346;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1552 <= 0;
  else
    g1552 <= g7347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1555 <= 0;
  else
    g1555 <= g7348;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1558 <= 0;
  else
    g1558 <= g7349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1561 <= 0;
  else
    g1561 <= g7350;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1564 <= 0;
  else
    g1564 <= g7351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1570 <= 0;
  else
    g1570 <= g4900;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1567 <= 0;
  else
    g1567 <= g7352;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1571 <= 0;
  else
    g1571 <= g7353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1574 <= 0;
  else
    g1574 <= g7354;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1577 <= 0;
  else
    g1577 <= g7355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1580 <= 0;
  else
    g1580 <= g7356;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1583 <= 0;
  else
    g1583 <= g7357;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1586 <= 0;
  else
    g1586 <= g7358;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1589 <= 0;
  else
    g1589 <= g7359;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1592 <= 0;
  else
    g1592 <= g7360;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1595 <= 0;
  else
    g1595 <= g7361;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1598 <= 0;
  else
    g1598 <= g7362;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1601 <= 0;
  else
    g1601 <= g7363;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1604 <= 0;
  else
    g1604 <= g7364;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1607 <= 0;
  else
    g1607 <= g7365;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1654 <= 0;
  else
    g1654 <= g10874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1657 <= 0;
  else
    g1657 <= g10875;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1660 <= 0;
  else
    g1660 <= g11033;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1663 <= 0;
  else
    g1663 <= g11034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1666 <= 0;
  else
    g1666 <= g11035;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1669 <= 0;
  else
    g1669 <= g11036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1672 <= 0;
  else
    g1672 <= g11037;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1675 <= 0;
  else
    g1675 <= g11038;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1678 <= 0;
  else
    g1678 <= g11039;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1681 <= 0;
  else
    g1681 <= g11040;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1684 <= 0;
  else
    g1684 <= g11041;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1687 <= 0;
  else
    g1687 <= g11042;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g546 <= 0;
  else
    g546 <= g11043;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g554 <= 0;
  else
    g554 <= g11047;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g557 <= 0;
  else
    g557 <= g11048;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g560 <= 0;
  else
    g560 <= g11049;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g563 <= 0;
  else
    g563 <= g11050;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g566 <= 0;
  else
    g566 <= g11051;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g569 <= 0;
  else
    g569 <= g10876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g572 <= 0;
  else
    g572 <= g10877;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g575 <= 0;
  else
    g575 <= g11052;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g549 <= 0;
  else
    g549 <= g11044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g552 <= 0;
  else
    g552 <= g11045;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g553 <= 0;
  else
    g553 <= g11046;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g23 <= 0;
  else
    g23 <= g3327;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g26 <= 0;
  else
    g26 <= g4885;
assign g2171 = ((~II5116));
assign g3491 = ((~g2669));
assign g2000 = ((~g810));
assign g10722 = (g10308)|(g10671);
assign II12647 = ((~g7711));
assign g6579 = ((~g5949));
assign g10241 = ((~g10192));
assign II13463 = ((~g8156));
assign II10924 = ((~g6736));
assign II12216 = ((~g2518))|((~II12214));
assign II14835 = (g9621)|(g9645)|(g9588);
assign g10306 = (g10214&g9082);
assign g4866 = (g231&g3946);
assign g10861 = (g5523)|(g10745);
assign g8600 = ((~g8475));
assign g3783 = ((~II7009));
assign g8117 = (g6236&g7886);
assign g8508 = (g8411&g7967);
assign g8487 = ((~g8350));
assign g6136 = ((~II9845));
assign g10300 = (g8892&g10220);
assign II4783 = ((~g873));
assign g7555 = ((~II11989));
assign g8588 = ((~II13831));
assign g11145 = (g315&g10927);
assign g7570 = ((~II12032));
assign g7881 = (g7612&g3810);
assign g7658 = ((~II12271));
assign g2776 = ((~II5866))|((~II5867));
assign II12226 = ((~g7066));
assign g9834 = (g9731&g9785);
assign g9621 = (g1179&g9125);
assign g6426 = ((~II10340));
assign g8278 = ((~II13206));
assign II10349 = ((~g6215));
assign II8711 = ((~g4530));
assign II7405 = ((~g3861));
assign g8946 = ((~II14295));
assign g10764 = (g10643&g4840);
assign g9700 = (g9358)|(g9667)|(II14827);
assign II5315 = ((~g1032))|((~g1027));
assign g8932 = ((~II14264))|((~II14265));
assign II7562 = ((~g3533))|((~g654));
assign g4960 = (g1403&g4682);
assign g9338 = ((~II14519));
assign g3221 = ((~g1834))|((~g2564));
assign g6045 = (g5541)|(g3989);
assign II5891 = ((~g750))|((~g2057));
assign g10695 = ((~II16366));
assign g11192 = (g5628&g11066);
assign g7246 = (g6465)|(g6003);
assign II7432 = ((~g3663));
assign g2039 = ((~g1781));
assign II16051 = ((~g837))|((~g10371));
assign g5845 = ((~g5320));
assign g2321 = ((~II5372))|((~II5373));
assign II10228 = ((~g6113));
assign II5095 = ((~g37));
assign g7440 = ((~II11836));
assign II5689 = (g1419&g1424&g1428&g1432);
assign g2662 = ((~g2014));
assign g7600 = ((~II12150));
assign II15871 = ((~g10358))|((~II15870));
assign g8801 = (g8742&g8729);
assign g7756 = ((~II12433));
assign g5119 = ((~II8514))|((~II8515));
assign g5099 = (g4821&g3829);
assign g7636 = ((~II12248));
assign II7441 = ((~g3473));
assign g10310 = ((~II15736));
assign g4097 = (g2677&g2989);
assign II10039 = ((~g5718));
assign g5778 = ((~II9368));
assign g8641 = (g8120)|(g8463);
assign g9606 = ((~g9125)&(~g9111)&(~g9173)&(~g9151));
assign g4157 = (g2713&g3055);
assign II16847 = ((~g10886));
assign g10947 = ((~II16708));
assign g8938 = (g8789)|(g8699);
assign g5913 = (g1041&g5320);
assign g8976 = ((~II14349));
assign g9901 = (g9893&g9392);
assign g6544 = (g1227&g6081);
assign g5589 = ((~II9001));
assign g10743 = (g10639&g4013);
assign gbuf10 = (g1736);
assign II11907 = ((~g6967))|((~g1474));
assign g4276 = ((~g4065)&(~g3261)&(~g2500));
assign g10950 = (g10788&g6355);
assign g2651 = ((~g2007));
assign g8941 = (g8796)|(g8706);
assign g7521 = ((~II11901));
assign g6358 = (g5841&g4441);
assign g10560 = (g10487&g4575);
assign g4897 = ((~II8256));
assign g3638 = ((~II6821));
assign II15542 = ((~g10065));
assign II11440 = ((~g6577));
assign II16332 = ((~g4997))|((~II16330));
assign g9830 = (g9725&g9785);
assign g11259 = (g11236)|(g11021);
assign g10668 = ((~g10563));
assign g9717 = (g1537&g9490);
assign II16161 = (g10479)|(g10478)|(g10477)|(g10475);
assign g8717 = ((~II14010));
assign g10877 = ((~II16601));
assign g6890 = (g6752&g6568);
assign g10732 = (g4358)|(g10661);
assign g9809 = ((~II14944));
assign gbuf3 = (g755);
assign II8562 = ((~g4227))|((~II8561));
assign g11545 = ((~g11519));
assign g10872 = ((~II16586));
assign II6631 = (g2707&g2713&g2719&g2765);
assign II17407 = ((~g11417));
assign g10783 = ((~II16479));
assign g2503 = ((~g1872));
assign g8106 = ((~g7950));
assign II7109 = ((~g2970));
assign g2135 = ((~II5064));
assign g10230 = (g8892&g10145);
assign II15187 = ((~g9968));
assign II5192 = ((~g55));
assign g6114 = ((~II9795));
assign II9804 = ((~g5417));
assign g11232 = (g11158)|(g11015);
assign II16550 = ((~g10726));
assign g6847 = ((~g6482));
assign g6818 = ((~II10864));
assign g10495 = (g10431&g3971);
assign g10685 = (g10608&g3863);
assign g5491 = (g1624&g4262);
assign g10882 = ((~II16616));
assign g8645 = (g8127)|(g8469);
assign II11436 = ((~g6488));
assign g4883 = (g248&g3946);
assign II17730 = ((~g11638));
assign g10186 = ((~II15536));
assign g6015 = (g5497)|(g3942);
assign g7136 = (g6050&g6704);
assign g4939 = ((~II8303));
assign g5726 = (g1601&g5167);
assign g2177 = ((~II5127))|((~II5128));
assign II16407 = ((~g10696));
assign II15281 = ((~g10025));
assign g9962 = (g9952&g9536);
assign g8885 = (g8841)|(g8754);
assign g6827 = (g219&g6596);
assign g8143 = ((~g8029));
assign g10778 = (g1027&g10729);
assign g5673 = ((~II9180));
assign g11650 = ((~II17752));
assign g8130 = (g1936&g7952);
assign II10507 = ((~g6221))|((~g786));
assign g5295 = ((~II8762))|((~II8763));
assign g6743 = (g4106&g6146);
assign g6101 = ((~II9762));
assign II6543 = ((~g3186));
assign II8256 = ((~g4711));
assign g11472 = ((~II17453));
assign g8123 = (g1918&g7946);
assign g7569 = ((~II12029));
assign g3748 = ((~g2971));
assign g6279 = ((~II10096));
assign g9109 = ((~II14452));
assign II12678 = ((~g7376));
assign g7942 = ((~g7395))|((~g6847))|((~g7380))|((~g7369));
assign g5318 = (g4401&g1857);
assign II11427 = ((~g6573));
assign g4919 = ((~II8290));
assign II11417 = ((~g6638));
assign g6594 = ((~II10560));
assign g8817 = (g7954)|(g8732);
assign II16540 = ((~g10722));
assign g8032 = (g7385&g7438);
assign II17243 = ((~g11396));
assign g9738 = (g9417)|(g9447)|(g9506);
assign g6155 = ((~g4974)&(~g2864));
assign g11584 = (g1318&g11542);
assign g7914 = ((~g7651));
assign g5602 = (g1624&g4535);
assign g1976 = ((~g643));
assign II4941 = ((~g396))|((~g324));
assign g9665 = (g1314&g9151);
assign g8704 = ((~g8667));
assign II9647 = ((~g5148));
assign II13544 = ((~g713))|((~g8259));
assign g2087 = ((~g225));
assign II15539 = ((~g10069));
assign II11773 = ((~g7257));
assign g6333 = (g197&g5904);
assign II13858 = ((~g8538))|((~II13857));
assign g2315 = (g1163)|(g1166)|(g1113)|(II5363);
assign g6108 = ((~II9779));
assign II8982 = ((~g4728));
assign g6389 = ((~II10289));
assign g10270 = ((~g10156));
assign g4899 = ((~II8262));
assign II12406 = ((~g7464));
assign g7264 = ((~II11501));
assign g3385 = ((~g3121));
assign g6364 = (g5851&g4454);
assign g8219 = ((~g7826));
assign g11575 = ((~g11561));
assign g3200 = ((~g1822))|((~g2061));
assign g5185 = ((~g4682));
assign g4459 = ((~II7820));
assign g9347 = ((~II14546));
assign g4717 = ((~g3829));
assign g8384 = (g8180&g3397);
assign g10217 = ((~II15589));
assign II15314 = ((~g10007));
assign g10025 = (II15224)|(II15225);
assign g4413 = ((~II7749));
assign g4127 = ((~II7276));
assign g10117 = ((~II15359));
assign g8804 = ((~II14133));
assign g5947 = ((~II9585));
assign II9259 = ((~g5301));
assign II5485 = ((~g1250))|((~II5484));
assign II13933 = ((~g8505));
assign g1982 = ((~g736));
assign II5391 = ((~g1101));
assign g10125 = ((~II15377));
assign II9893 = ((~g5557));
assign g7818 = (g1878&g7479);
assign g5935 = ((~II9558))|((~II9559));
assign g10134 = ((~II15400));
assign g6086 = ((~II9737));
assign g7297 = (g7132)|(g6323);
assign g11266 = (g11190)|(g11028);
assign g11331 = (g11272)|(g11171);
assign g5258 = (g700&g4756);
assign II5500 = ((~g1255))|((~g1007));
assign g2941 = ((~II6118));
assign g3990 = ((~g3121));
assign g2727 = ((~g2022));
assign g10894 = ((~II16644));
assign g2340 = ((~g1918));
assign g9451 = ((~II14642));
assign g2054 = ((~g1864));
assign g7132 = (g6048&g6702);
assign II16766 = ((~g10892));
assign g7797 = ((~II12556));
assign II13714 = ((~g8351));
assign g1989 = ((~g770));
assign g9709 = (g1524&g9490);
assign g9360 = ((~II14579));
assign g8210 = (g7466)|(g7995);
assign g6822 = (g231&g6596);
assign II8831 = ((~g4480));
assign g7409 = (g4976&g632&g6858);
assign g10400 = ((~g10348));
assign II15060 = ((~g9696));
assign g8044 = (g7598&g5919);
assign II5792 = ((~g2080));
assign II7665 = ((~g3732));
assign II6901 = ((~g2818));
assign g11284 = ((~g11208));
assign g2984 = (g2528)|(g2522);
assign II14449 = ((~g8973));
assign g8137 = ((~II13010));
assign g5512 = (g1660&g4281);
assign g10405 = (g10297)|(g9530);
assign g4461 = ((~g3829));
assign g4168 = ((~II7322))|((~II7323));
assign g6488 = ((~g6027))|((~g6019));
assign II14271 = ((~g8840))|((~II14270));
assign g4720 = (g1023&g3914);
assign g7588 = ((~II12093))|((~II12094));
assign g6150 = ((~II9869));
assign II6643 = ((~g3008));
assign g7537 = ((~II11947));
assign g9868 = (g1555&g9812);
assign g6662 = (g366&g6220);
assign g5489 = (g4287&g3521);
assign g6269 = ((~II10066));
assign g3109 = ((~g2482));
assign g9582 = (g2725&g9173);
assign g2181 = ((~II5142));
assign g4999 = (g1499&g4640);
assign g11032 = (g416&g10974);
assign II8333 = ((~g4456));
assign g7962 = (g7730&g6712);
assign g2328 = ((~g1882));
assign g9696 = (g281&g9432);
assign g5305 = ((~g4378));
assign II9341 = ((~g5013));
assign g9357 = (g962&g9223);
assign II7303 = ((~g3262));
assign II13962 = ((~g8451));
assign II13341 = ((~g8210));
assign g9914 = (g9851)|(g9692);
assign g8461 = (g8298&g7403);
assign g2157 = ((~g1703));
assign II17337 = ((~g11363));
assign g2014 = ((~g1104));
assign g11633 = ((~II17713));
assign II12085 = ((~g6980))|((~g1470));
assign g6536 = ((~II10456));
assign g11169 = (g530&g11112);
assign g9271 = (g6681&g8949);
assign g8556 = (g8412&g8029);
assign g10201 = ((~g10175));
assign g4064 = (g1759&g2799);
assign g8250 = (g2771&g7907);
assign g8982 = ((~II14367));
assign g3807 = (g3003&g3062);
assign g10453 = (g10437&g3395);
assign II14506 = ((~g8923));
assign g6900 = (g6787)|(g6246);
assign g2669 = ((~g2015));
assign g5074 = (g1771&g4587);
assign II5085 = (g1490&g1494&g1504&g1508);
assign g3213 = ((~II6388));
assign II5459 = ((~g1240))|((~g1003));
assign II10042 = ((~g5723));
assign g9683 = (g9454)|(g9292)|(g9274);
assign g11344 = ((~II17155));
assign g7681 = ((~g7148));
assign g2733 = ((~II5795));
assign II11330 = ((~g6571));
assign II14855 = (g9583)|(g9593)|(g9601)|(g9596);
assign II6861 = ((~g2942));
assign II9279 = ((~g5314));
assign g2462 = ((~II5555));
assign II17563 = ((~g11492));
assign g2246 = ((~g1810));
assign g11506 = ((~II17537));
assign g11484 = (g6639)|(g11461);
assign g4777 = ((~g3992));
assign II6414 = ((~g2342));
assign II9992 = ((~g5633));
assign II7577 = ((~g4124));
assign g5525 = (g1721&g4292);
assign g11006 = (g5125&g10827);
assign g6654 = (g363&g6214);
assign g10328 = (g10252&g3307);
assign g5815 = ((~II9421));
assign g3991 = (g1738&g2774);
assign II15858 = ((~g10336));
assign g4637 = ((~II8039));
assign g7364 = ((~II11740));
assign II10048 = ((~g5734));
assign g2025 = ((~g1696));
assign g11613 = (g11600)|(g11591);
assign II13430 = ((~g8241));
assign g9825 = ((~II14976));
assign II7487 = ((~g3371));
assign g4285 = ((~g3688));
assign II11524 = ((~g6593));
assign g7316 = ((~II11596));
assign g5274 = ((~II8729))|((~II8730));
assign g2614 = ((~g1994));
assign II15042 = (g7853)|(g9686)|(g9624)|(g9785);
assign g6961 = ((~II11115));
assign g10527 = ((~g10462));
assign g7339 = ((~II11665));
assign g2211 = ((~g153));
assign g5210 = ((~II8631));
assign g11045 = ((~II16796));
assign g8206 = (g7459)|(g8007);
assign g6225 = (g566&g5082);
assign g3051 = ((~g2135));
assign II9680 = ((~g5194));
assign g5820 = (g5595)|(g4834);
assign II16203 = ((~g10454));
assign g7747 = ((~II12406));
assign g10279 = ((~g10158));
assign g11163 = ((~II16920));
assign g4468 = ((~II7837));
assign g3066 = ((~g2135));
assign II6225 = ((~g2544))|((~II6224));
assign g5268 = (g1098&g4769);
assign g6416 = (g3497&g5774);
assign g5038 = (g4878)|(g4884);
assign g8159 = (g7895)|(g6886);
assign g3463 = ((~g3256));
assign g7896 = ((~II12678));
assign II16360 = ((~g10590));
assign II14315 = ((~g8815));
assign g4508 = ((~g3946));
assign g11342 = ((~II17149));
assign II10801 = ((~g6536));
assign g7386 = ((~II11767));
assign g10373 = ((~g10346)&(~g3463));
assign g8293 = ((~II13233));
assign g7449 = (g6868&g4355);
assign II15778 = ((~g10255));
assign II5237 = ((~g1107));
assign II15311 = ((~g10013));
assign II12193 = ((~g7270));
assign II16979 = ((~g11088));
assign g7024 = ((~II11169));
assign g10969 = (g3625&g10809);
assign II9639 = ((~g5126));
assign g6176 = ((~II9905));
assign II9020 = ((~g4773));
assign g4972 = (g1436&g4682);
assign II10398 = ((~g5820));
assign II13523 = ((~g8249))|((~II13521));
assign II10834 = ((~g6715));
assign g6909 = (g6346)|(g5684);
assign g11081 = ((~II16856));
assign II5064 = ((~g1690));
assign g2683 = ((~g2037));
assign II5667 = ((~g566));
assign g10762 = (g10635&g4840);
assign g11080 = ((~II16853));
assign II6742 = ((~g3326));
assign g3398 = ((~g2896));
assign g7787 = ((~II12526));
assign g4267 = ((~g3800)&(~g2593)&(~g2586)&(~g2579));
assign II11034 = ((~g6629));
assign g3144 = ((~g2462));
assign II5510 = ((~g588));
assign g10972 = ((~II16717));
assign II13230 = ((~g8244));
assign g7143 = (g6619)|(g6039);
assign g10332 = ((~II15782));
assign II12550 = ((~g7675));
assign g10770 = (g5525)|(g10682);
assign g6884 = (g5569&g6564);
assign II16679 = ((~g10784));
assign II15962 = ((~g10405));
assign g3475 = ((~g3056));
assign g11491 = ((~II17493))|((~II17494));
assign g7147 = ((~II11394));
assign g6049 = (g5254)|(g3718);
assign II15861 = ((~g10339));
assign g10007 = (II15209)|(II15210);
assign II6156 = ((~g2119));
assign II7877 = ((~g810))|((~II7875));
assign g7593 = ((~II12114))|((~II12115));
assign g11550 = ((~II17591));
assign g9111 = (g8965&g6674);
assign g7676 = ((~II12303));
assign g4732 = (g391&g3372);
assign II15256 = ((~g9984))|((~g9980));
assign g10854 = ((~g10708));
assign II13738 = ((~g8295));
assign g10333 = (g10262&g3307);
assign II17453 = ((~g11451));
assign II11992 = ((~g7058));
assign g5894 = ((~g5361));
assign g10384 = ((~II15871))|((~II15872));
assign g2334 = ((~II5388));
assign g11260 = (g11237)|(g11022);
assign II13695 = ((~g8363));
assign g10616 = ((~II16289));
assign g2990 = (g2061&g2557&g1814);
assign II10958 = ((~g6559));
assign g3697 = ((~II6856));
assign II10546 = ((~g5914));
assign g10543 = ((~II16196));
assign g7734 = (g6944&g3880);
assign II17225 = ((~g11298));
assign II6031 = ((~g2209));
assign II10598 = ((~g5874));
assign g7761 = ((~II12448));
assign g6252 = ((~II10015));
assign II13831 = ((~g8560));
assign g4435 = ((~g3914));
assign II10421 = ((~g5826));
assign g8891 = ((~II14239));
assign II5441 = ((~g919));
assign g5766 = ((~II9346));
assign II13083 = ((~g7921));
assign g4283 = (g4059)|(g4063);
assign g10165 = ((~II15491));
assign II9240 = ((~g5069));
assign g4824 = (g774&g4099);
assign g7075 = (g5104)|(g6530);
assign g2864 = ((~g2298));
assign II10168 = ((~g5982));
assign g10545 = ((~II16200));
assign g7049 = ((~II11228));
assign g11108 = ((~g10974));
assign g8640 = ((~g8512));
assign g6569 = ((~II10499));
assign g9919 = ((~II15114));
assign g5624 = ((~II9056));
assign g2771 = ((~II5854));
assign g8844 = (g8609&g8709);
assign g8837 = (g8646&g8697);
assign g8664 = ((~II13949));
assign g7137 = (g5590&g6361);
assign II9550 = ((~g5030));
assign g2482 = ((~II5565));
assign g11022 = (g444&g10974);
assign II6454 = ((~g2368));
assign g11224 = (g968&g11056);
assign g7390 = ((~g6847));
assign II5662 = ((~g563));
assign g4219 = ((~g3635));
assign g4790 = ((~g3337));
assign g9876 = ((~g9522)&(~g9536)&(~g9576)&(~II15039));
assign II13125 = ((~g7975));
assign g3517 = ((~II6702));
assign II15088 = ((~g9832));
assign II11397 = ((~g6713));
assign g9448 = ((~g9091));
assign II11149 = ((~g6468));
assign g8565 = ((~II13788));
assign II15782 = ((~g10259));
assign g3585 = ((~II6747))|((~II6748));
assign II16708 = ((~g10822));
assign g7307 = ((~II11569));
assign g10140 = ((~II15418));
assign g11324 = (g11271)|(g11164);
assign II5373 = ((~g976))|((~II5371));
assign g4170 = ((~g3328));
assign II5632 = ((~g932));
assign g6804 = ((~II10822));
assign g10729 = ((~g10630));
assign g2253 = ((~g100));
assign g7908 = ((~g7454));
assign g3375 = ((~II6569));
assign II11176 = ((~g6501));
assign g3874 = ((~g2920));
assign g11196 = (g4912&g11068);
assign II6598 = ((~g2623));
assign II8671 = ((~g814))|((~II8669));
assign II15403 = ((~g10069));
assign II9352 = ((~g4944));
assign g6899 = (g6463)|(g5471);
assign g10750 = (g10687&g3586);
assign II9938 = ((~g5478));
assign g10692 = ((~II16363));
assign g5010 = (g1458&g4640);
assign g5650 = ((~II9111));
assign II10816 = ((~g6406));
assign g6670 = ((~II10633));
assign g6465 = (g5825)|(g5041);
assign II17149 = ((~g11306));
assign g5251 = ((~g4640));
assign g10092 = ((~II15323));
assign g10043 = ((~II15257))|((~II15258));
assign II10090 = ((~g5767));
assign g5405 = (g4476)|(g3440);
assign g10503 = (g10388&g2135);
assign g4678 = ((~g3546));
assign g5630 = ((~II9068));
assign g7709 = (g6856&g4333);
assign g3631 = ((~II6793))|((~II6794));
assign g3726 = ((~II6898));
assign g7950 = ((~g7395))|((~g7390))|((~g7380))|((~g7273));
assign II5403 = ((~g636));
assign II12613 = ((~g7525));
assign II16239 = ((~g10525));
assign II15085 = ((~g9720));
assign g11295 = (g5475&g11239);
assign II12478 = ((~g7560));
assign g6260 = ((~II10039));
assign II13272 = ((~g1918))|((~g8158));
assign II7288 = ((~g2873));
assign g6679 = (g4631&g6074&g2733);
assign II14094 = ((~g8700));
assign g2373 = ((~g471));
assign II17461 = ((~g11448))|((~II17459));
assign g6064 = (g5398&g2230);
assign g2918 = (g2411&g1672);
assign g2959 = ((~II6167))|((~II6168));
assign II16613 = ((~g10794));
assign g4873 = ((~g3292)&(~g2593)&(~g2586)&(~g3776));
assign II14228 = ((~g8797));
assign g7330 = ((~II11638));
assign g3945 = ((~II7096));
assign g4596 = ((~II8007));
assign g4613 = ((~g3077)&(~g3491)&(~g2662)&(~g2655));
assign g6771 = (g263&g5866);
assign g11616 = ((~II17666));
assign g11241 = ((~g11112));
assign g8131 = ((~g8020));
assign g7610 = ((~II12180));
assign g10265 = ((~g10143));
assign g8446 = ((~II13636));
assign g8781 = ((~II14080));
assign g9426 = ((~g9052)&(~g9030));
assign g6553 = ((~II10477));
assign g10794 = ((~II16496));
assign II13239 = ((~g8266));
assign g4048 = (g1750&g2790);
assign II14522 = ((~g9108));
assign II8869 = ((~g4421));
assign g8426 = ((~II13592));
assign II14263 = ((~g8843))|((~g1814));
assign II12989 = ((~g8043));
assign g11304 = (g5520&g11245);
assign II8154 = ((~g3636));
assign g5882 = (g5592&g3829);
assign g4840 = ((~II8199));
assign g5486 = ((~g4395));
assign II11058 = ((~g6641));
assign II6085 = ((~g2234));
assign II8303 = ((~g4784));
assign g2647 = ((~g1993));
assign II11228 = ((~g6471));
assign II13723 = ((~g8359));
assign g8152 = ((~II13043));
assign II8178 = ((~g3685))|((~g1786));
assign g3118 = ((~g2521)&(~g2514));
assign g9566 = (g9052)|(g9030);
assign II9559 = ((~g782))|((~II9557));
assign g8501 = ((~g3760))|((~g8366));
assign g3721 = ((~II6891));
assign g2406 = ((~g1365));
assign g5747 = ((~II9317));
assign g10463 = ((~II15980));
assign g8335 = ((~II13385));
assign g7268 = ((~II11505));
assign II6996 = ((~g2904));
assign g9366 = (g1311&g9173);
assign g6308 = ((~II10183));
assign g7656 = ((~II12265));
assign g11230 = (g471&g11062);
assign g8434 = (g8400)|(g8074);
assign II12832 = ((~g7681));
assign g2203 = ((~g677));
assign II7701 = ((~g3513));
assign II8320 = ((~g4452));
assign II8240 = ((~g4380));
assign g2541 = ((~II5658));
assign II6488 = ((~g2306))|((~II6487));
assign g1998 = ((~g802));
assign g3228 = ((~II6409));
assign g3903 = ((~II7070));
assign g2354 = ((~g1515))|((~g1520));
assign g5864 = ((~II9483));
assign II10702 = ((~g6071));
assign II8631 = ((~g4425));
assign g8962 = (g8089&g6368&g8828);
assign II16095 = ((~g10401));
assign II15729 = ((~g10254));
assign g7070 = ((~II11289));
assign g3076 = ((~II6282));
assign II5135 = ((~g521))|((~g525));
assign II6406 = ((~g2339));
assign g7894 = (g7617&g3816);
assign II16629 = ((~g10860));
assign g5395 = ((~II8831));
assign II13589 = ((~g8361));
assign II8436 = ((~g4462));
assign g5689 = ((~II9216));
assign g7191 = (g6343&g4323);
assign g9716 = (g1534&g9490);
assign g11046 = ((~II16799));
assign II12535 = ((~g7656));
assign II7354 = ((~g4066));
assign g2832 = ((~II5946));
assign II13669 = ((~g8294));
assign II7633 = ((~g3474));
assign II17513 = ((~g11482));
assign II8590 = ((~g4251))|((~II8589));
assign II13822 = ((~g8488));
assign g4054 = (g1753&g2793);
assign II11106 = ((~g6667));
assign II12143 = ((~g7089))|((~g158));
assign g2964 = ((~II6193));
assign g10348 = (g10272&g3705);
assign II10666 = ((~g6042));
assign g10177 = ((~II15523));
assign g11586 = (g1324&g11545);
assign g10575 = ((~g10523));
assign II9199 = ((~g4935));
assign g7213 = ((~II11447));
assign g10175 = ((~II15517));
assign g8768 = (g8623&g5151);
assign g5984 = ((~II9602));
assign g7358 = ((~II11722));
assign g6094 = ((~II9749));
assign II5015 = ((~g1011))|((~II5013));
assign g9124 = (g8881&g4802);
assign g9262 = ((~II14473));
assign g4213 = ((~II7456));
assign g6924 = (g6362)|(g4261);
assign II7779 = ((~g3774));
assign g6070 = (g1050&g5320);
assign g11222 = (g965&g11055);
assign g4730 = ((~g3546));
assign g3459 = ((~II6661));
assign g3291 = ((~g2161));
assign II9008 = ((~g1791))|((~II9006));
assign g9595 = (g901&g9205);
assign g7603 = ((~II12159));
assign g4094 = ((~g2744));
assign g7884 = (g7457&g7022);
assign II12127 = ((~g7103))|((~II12126));
assign II8513 = ((~g4873))|((~g3513));
assign II14236 = ((~g8802));
assign g6541 = (g5788)|(g5009);
assign II5588 = ((~g1203));
assign g6995 = ((~g6482));
assign g3435 = (g2945)|(g2950);
assign II12916 = ((~g7849));
assign II13096 = ((~g7925));
assign g10880 = ((~II16610));
assign g5693 = ((~II9224));
assign g2222 = ((~g158));
assign g11311 = ((~II17100));
assign II6439 = ((~g2352));
assign g2891 = ((~II6055));
assign g7972 = ((~II12770));
assign g10204 = ((~g10174));
assign g2369 = ((~g617));
assign g7011 = ((~g6503));
assign II11713 = ((~g7023));
assign g6970 = ((~II11122));
assign II5943 = ((~g2233));
assign g8418 = ((~II13568));
assign II4906 = ((~g119));
assign g10667 = (g10576&g9427);
assign II5989 = ((~g2252));
assign II11980 = ((~g6957))|((~g1482));
assign g6248 = ((~II10003));
assign g4307 = ((~g4013));
assign g2607 = ((~II5722));
assign g8883 = (g8838)|(g8753);
assign g10440 = ((~g10360))|((~g6037));
assign g10507 = ((~g10434))|((~g5859));
assign g4343 = (g345&g3586);
assign II16802 = ((~g10902));
assign II13391 = ((~g8178));
assign g11237 = (g5472&g11109);
assign II9001 = ((~g4762));
assign g8362 = ((~II13466));
assign g5875 = ((~g5361));
assign g10194 = ((~g10062));
assign g10536 = ((~II16175));
assign g11248 = (g976&g11071);
assign g11070 = (g2008&g10913);
assign II14613 = ((~g9204))|((~II14612));
assign g7926 = (g7435)|(g6892);
assign II12773 = ((~g7581));
assign g5514 = (g1941&g4284);
assign g8069 = (g673&g7826);
assign g11557 = (g2707&g11519);
assign g7227 = ((~II11467));
assign g9512 = (g9151)|(g9125);
assign g2274 = ((~II5324))|((~II5325));
assign II6178 = ((~g197))|((~II6176));
assign II12239 = ((~g7073));
assign II9162 = ((~g5035));
assign II17185 = ((~g11311));
assign g2548 = ((~II5667));
assign g5026 = (g1453&g4640);
assign g11306 = (g11216)|(g11095);
assign g11062 = ((~g10937));
assign g5682 = ((~II9199));
assign II11405 = ((~g6627));
assign g4395 = ((~II7732));
assign g8187 = (g7542)|(g7998);
assign g8846 = (g8615&g8712);
assign g3685 = (g1781&g2981);
assign II15356 = ((~g10013));
assign g2213 = ((~g1110));
assign II5734 = ((~g2097));
assign g5547 = (g1733&g4326);
assign II12770 = ((~g7638));
assign g10339 = (g10232)|(g9556);
assign II8449 = ((~g4469));
assign II6958 = ((~g2872));
assign g3343 = ((~g2779));
assign II6528 = ((~g3274));
assign II10633 = ((~g6015));
assign g11155 = ((~g10950));
assign II9302 = ((~g5576));
assign g5446 = ((~II8877));
assign g6309 = ((~II10186));
assign g9758 = ((~g9454)&(~g9274)&(~g9292));
assign g10902 = ((~II16660));
assign g11033 = ((~II16760));
assign g3068 = ((~g2303));
assign g10466 = ((~II15989));
assign g7377 = ((~II11759));
assign g2858 = ((~II5992));
assign g9029 = ((~II14424));
assign g7791 = ((~II12538));
assign g6395 = ((~II10293));
assign II15412 = ((~g10075));
assign g4115 = (g2689&g3009);
assign g10188 = ((~II15542));
assign II17402 = ((~g11416))|((~II17400));
assign g7531 = ((~II11929));
assign g3332 = ((~II6513));
assign g3396 = (g213&g3228);
assign II11315 = ((~g6644));
assign g5477 = (g1887&g4241);
assign g3095 = ((~g2482));
assign g10365 = (g10319&g2135);
assign g5062 = ((~g4840));
assign g3437 = ((~II6654));
assign g10624 = (g10545&g4544);
assign g8788 = ((~II14097));
assign g11630 = ((~II17704));
assign II10563 = ((~g6043));
assign g7185 = (g1887&g6724);
assign g5149 = ((~II8551));
assign g7538 = ((~II11950));
assign II5231 = ((~g148))|((~II5229));
assign g5540 = (g1727&g4315);
assign g5888 = ((~g5102));
assign g3911 = ((~g3015));
assign II11132 = ((~g6451));
assign g3760 = ((~g3003));
assign g4321 = ((~g3863));
assign g2239 = ((~II5240));
assign g6186 = (g546&g5042);
assign g11363 = ((~II17188));
assign g5277 = ((~g3734))|((~g4538));
assign II13571 = ((~g8355));
assign II12583 = ((~g7546));
assign g3767 = ((~II6976));
assign g8727 = ((~g8592));
assign II11786 = ((~g7246));
assign g8557 = (g8415&g8033);
assign g7022 = ((~g6389));
assign II7790 = ((~g3782));
assign g4179 = ((~II7354));
assign g5197 = ((~II8611));
assign g5217 = ((~II8641))|((~II8642));
assign g2111 = ((~II5006))|((~II5007));
assign II10736 = ((~g6104));
assign g7935 = (g2821&g7454);
assign g4601 = ((~g3077)&(~g2669)&(~g2662)&(~g3479));
assign g6200 = ((~II9935));
assign g3792 = ((~II7017));
assign g3383 = (g186&g3228);
assign II6167 = ((~g2236))|((~II6166));
assign g8402 = ((~II13505))|((~II13506));
assign g7678 = ((~II12307));
assign g10594 = ((~g10480)&(~g10521));
assign II12020 = ((~g7119))|((~II12019));
assign g9751 = (g9515)|(g9510);
assign II9795 = ((~g5404));
assign g9385 = (g1324&g9151);
assign II17504 = ((~g11475))|((~II17503));
assign g4669 = ((~g4013));
assign II10519 = ((~g6231))|((~g822));
assign g9936 = (g9915&g9624);
assign g3429 = (g231&g3228);
assign g7458 = ((~g7123));
assign g6588 = ((~II10546));
assign g2079 = ((~II4891));
assign II5080 = ((~g36));
assign II12652 = ((~g7458));
assign g3327 = ((~II6498));
assign II17307 = ((~g11377))|((~II17305));
assign II9872 = ((~g5557));
assign g7810 = ((~II12595));
assign II7225 = ((~g1781))|((~II7223));
assign II6825 = ((~g3281))|((~g770));
assign II14439 = ((~g8969));
assign g7056 = ((~II11249));
assign g4221 = ((~g3914));
assign II16510 = ((~g10712));
assign g10911 = ((~II16685));
assign g6524 = (g5746)|(g4996);
assign II5120 = ((~g622));
assign g6196 = ((~g5446));
assign II9869 = ((~g5405));
assign II6894 = ((~g2813));
assign g10581 = (g10531&g9453);
assign g6941 = ((~g6503));
assign g6077 = ((~II9720));
assign II16871 = ((~g10973));
assign g9052 = (g8936&g7192);
assign II4891 = ((~g582));
assign g11455 = (g11435&g5446);
assign g9667 = ((~g9125)&(~g9111)&(~g9173)&(~g9151));
assign g6685 = ((~II10648));
assign g9956 = (g9948)|(g9942)|(g9815);
assign g9766 = ((~g9432));
assign II10308 = ((~g6003));
assign g3405 = ((~g3144));
assign g2306 = (g1223&g1218);
assign g8072 = (g700&g7826);
assign II15127 = ((~g9919));
assign g6392 = ((~g5859)&(~g5938));
assign g10438 = ((~g10356)&(~g3566));
assign g5231 = ((~g4640));
assign II15275 = ((~g9994));
assign II7393 = ((~g4096));
assign g4309 = (g4069)|(g4079);
assign g2509 = ((~II5588));
assign g5995 = (g5097)|(g5099);
assign II6971 = ((~g2882));
assign g5782 = (g1558&g5223);
assign II9786 = ((~g5396));
assign g8985 = ((~II14376));
assign II14087 = ((~g8770));
assign g10599 = (g10534&g4365);
assign g8550 = (g8402&g8011);
assign g10475 = ((~II16031))|((~II16032));
assign g4237 = ((~g4013));
assign g7937 = (g7606&g4013);
assign II6061 = ((~g2246));
assign II12809 = ((~g7686));
assign g2571 = ((~g1822));
assign II17662 = ((~g11602));
assign g3626 = ((~II6778))|((~II6779));
assign II5646 = ((~g940));
assign g9257 = (g6689&g8964);
assign g6530 = (g6207&g3829);
assign II6124 = ((~g2215))|((~g1419));
assign g8953 = ((~II14312));
assign II8651 = ((~g4824))|((~II8650));
assign g5069 = ((~g4368));
assign g2456 = ((~g1397));
assign II7360 = ((~g4081));
assign g8978 = ((~II14355));
assign g4226 = ((~g3698));
assign g8926 = (g8848)|(g8764);
assign II16277 = ((~g10536));
assign II12786 = ((~g7622));
assign II11674 = ((~g7051));
assign II6118 = ((~g2248));
assign II9232 = ((~g4944));
assign g2043 = ((~g1801));
assign II12526 = ((~g7648));
assign g4411 = ((~II7743));
assign g4755 = ((~g3440));
assign II8311 = ((~g4794));
assign g10699 = ((~II16376));
assign g9533 = ((~II14684));
assign g6322 = (g1275&g5949);
assign g10935 = ((~g10827));
assign g6207 = ((~II9947))|((~II9948));
assign g11013 = (g5209&g10827);
assign g9598 = (g2086&g9274);
assign II17543 = ((~g11499));
assign II14884 = ((~g9454));
assign II13406 = ((~g8179));
assign g3415 = ((~g3121));
assign II7863 = ((~g4099))|((~g774));
assign g8163 = (g7960&g3737);
assign g10019 = (II15219)|(II15220);
assign II15389 = ((~g10110));
assign g7702 = ((~g7079));
assign g3120 = (II6350)|(II6351);
assign II10021 = ((~g5692));
assign g8167 = (g5253&g7853);
assign II16220 = ((~g10502));
assign II13682 = ((~g8310));
assign g2554 = ((~II5672));
assign g8341 = ((~II13403));
assign g6698 = ((~II10671));
assign g11377 = ((~II17202));
assign II6385 = ((~g2260));
assign g10515 = (g10505&g10469&II16142);
assign g7752 = ((~II12421));
assign II16331 = ((~g10616))|((~II16330));
assign g10483 = ((~II16087))|((~II16088));
assign g9742 = (g9173)|(g9528);
assign II6025 = ((~g2259));
assign g10427 = ((~g10296)&(~g4620));
assign g4196 = ((~II7405));
assign g10649 = (g10626)|(g7741);
assign II9126 = ((~g4891));
assign g4457 = ((~g3829));
assign g11167 = (g538&g11112);
assign g9351 = ((~II14558));
assign II11596 = ((~g6831));
assign II9754 = ((~g5271));
assign g5574 = ((~g4300));
assign g11388 = ((~II17213));
assign II6665 = ((~g2792))|((~II6664));
assign II10678 = ((~g5777));
assign g10806 = ((~II16518));
assign g5202 = ((~g4640));
assign g10524 = ((~g10458));
assign g7201 = ((~II11427));
assign g11400 = ((~II17243));
assign II12508 = ((~g7731));
assign g6799 = ((~II10807));
assign g10255 = ((~g10139));
assign g5526 = (g1950&g4294);
assign g6435 = ((~II10355));
assign g11431 = ((~II17344));
assign II12344 = ((~g7062));
assign II9915 = ((~g5304));
assign g7906 = ((~II12694));
assign g7544 = ((~II11964));
assign g8710 = (g7607&g8595);
assign II11112 = ((~g6445));
assign g10396 = ((~II15907))|((~II15908));
assign II5652 = ((~g554));
assign g8081 = ((~g8000));
assign II16058 = ((~g841))|((~g10372));
assign II10015 = ((~g5641));
assign g10727 = (g4969)|(g10638);
assign II13869 = ((~g1403))|((~II13867));
assign g4513 = ((~g3546));
assign g2411 = ((~II5494));
assign g11515 = ((~g11490));
assign g7726 = ((~II12363));
assign II6467 = ((~g23))|((~g2479));
assign g9643 = (g950&g9223);
assign g6858 = ((~II10931))|((~II10932));
assign g11316 = (g11226)|(g11103);
assign g6302 = ((~II10165));
assign g8052 = (g7573&g5128);
assign g8005 = (g7510&g6871);
assign g4388 = ((~II7719));
assign g4312 = ((~g4144));
assign g6706 = ((~II10685));
assign II11238 = ((~g6543));
assign g11051 = ((~II16814));
assign g9950 = (g9901)|(g9898)|(g9779);
assign g10287 = ((~g10275)&(~g3463));
assign II17198 = ((~g11319));
assign II10120 = ((~g6248));
assign g10321 = ((~II15759));
assign II6173 = ((~g2125));
assign g11651 = ((~II17755));
assign II7163 = ((~g2643));
assign g10679 = ((~g10584));
assign II16190 = ((~g10493));
assign g8354 = ((~II13442));
assign II7964 = ((~g3433));
assign g5178 = (g2047&g4401&g4104);
assign II17340 = ((~g11366));
assign g5125 = ((~II8528))|((~II8529));
assign II8136 = ((~g4144));
assign II17282 = ((~g11360))|((~II17281));
assign g11188 = (g5604&g11063);
assign g4206 = ((~II7435));
assign g9525 = ((~g9257));
assign II10003 = ((~g4908));
assign II8763 = ((~g1129))|((~II8761));
assign g7320 = ((~II11608));
assign g9659 = (g956&g9223);
assign g4997 = (g4581)|(g4584);
assign g4161 = (g2719&g3060);
assign g5228 = (g1086&g4734);
assign g6660 = ((~II10623));
assign g2260 = ((~II5296))|((~II5297));
assign II9816 = ((~g5576));
assign g10229 = ((~II15608))|((~II15609));
assign g11541 = ((~g11519));
assign g6472 = (g5853&g1936);
assign II9576 = ((~g818))|((~II9574));
assign II12466 = ((~g7585));
assign g6764 = ((~g5987));
assign g2379 = (g744&g743);
assign g6747 = (g2214&g5897);
assign g5537 = (g4143&g4299);
assign II8414 = ((~g4293));
assign g3044 = ((~II6256));
assign g6314 = ((~II10201));
assign II17152 = ((~g11308));
assign g10630 = ((~II16311));
assign g9672 = ((~II14805));
assign g6368 = ((~g5987));
assign g2475 = ((~g192));
assign II8544 = ((~g4218))|((~II8543));
assign II6209 = ((~g802))|((~II6207));
assign g3262 = ((~II6432));
assign II11841 = ((~g7226));
assign g5120 = ((~II8520));
assign II11024 = ((~g6399));
assign g4482 = ((~II7864))|((~II7865));
assign II17176 = ((~g11286));
assign g4948 = ((~II8315));
assign g4901 = ((~II8268));
assign g11621 = ((~II17681));
assign g4764 = (g411&g3404);
assign g4559 = (g2034&g3829);
assign g7053 = ((~II11238));
assign g8327 = ((~g8164));
assign g4067 = ((~II7194));
assign g10739 = (g10676&g3368);
assign g8994 = (g8110&g6778&g8925);
assign II9498 = ((~g5081));
assign II13840 = ((~g8488));
assign II16775 = ((~g10889));
assign g11102 = (g861&g10950);
assign g10308 = (g10217&g9085);
assign g10512 = (g10395&g2135);
assign g10675 = ((~g10574));
assign g4503 = (g654&g3943);
assign II12463 = ((~g7579));
assign II10129 = ((~g5688));
assign g10294 = ((~II15704));
assign II11737 = ((~g7027));
assign II7825 = ((~g3414));
assign II5789 = ((~g2162));
assign gbuf5 = (g875);
assign II5171 = ((~g1419));
assign g6841 = (g1400&g6596);
assign g7066 = ((~II11275));
assign g5003 = (g1466&g4640);
assign g9100 = ((~g8892));
assign g6871 = ((~g6724));
assign II11858 = ((~g6888));
assign II10384 = ((~g5842));
assign II13078 = ((~g7963))|((~II13076));
assign g3817 = ((~II7043));
assign g5804 = (g1546&g5261);
assign g6617 = ((~g6019));
assign g10447 = ((~g10363))|((~g5360));
assign II15989 = ((~g10417));
assign g5787 = ((~II9383));
assign II6277 = ((~g1206));
assign g10639 = (g10623)|(g7734);
assign g7803 = ((~II12574));
assign g9894 = ((~II15085));
assign II5979 = ((~g2543));
assign II7402 = ((~g4121));
assign g9776 = ((~g9392)&(~g9367));
assign II17531 = ((~g11488));
assign II11286 = ((~g6551));
assign g10926 = ((~g10827));
assign g4095 = ((~II7233));
assign II15359 = ((~g10019));
assign II10132 = ((~g5696));
assign g6736 = ((~II10739));
assign g10301 = (g8892&g10223);
assign II15365 = ((~g10025));
assign g4181 = ((~II7360));
assign g4240 = ((~g3664));
assign g8288 = (g8119)|(g7825);
assign g2083 = ((~g139));
assign g3257 = (g378&g2496);
assign g8471 = ((~II13660))|((~II13661));
assign g2907 = ((~II6074));
assign g6255 = ((~II10024));
assign g9316 = (g8877&g5708);
assign II6793 = ((~g2959))|((~II6792));
assign g11438 = ((~II17365));
assign g6792 = (g290&g5881);
assign g9421 = ((~g9052)&(~g9030));
assign II17324 = ((~g11347));
assign II8796 = ((~g4672))|((~II8795));
assign g11207 = ((~II16982));
assign g5170 = (g1811&g4680);
assign g10730 = ((~II16407));
assign II11563 = ((~g6819));
assign g10825 = ((~II16537));
assign g9602 = (g2650&g9010);
assign g6217 = (g563&g5073);
assign g11336 = (g11281)|(g11176);
assign g11069 = ((~g10974));
assign g5847 = (g5626)|(g4877);
assign II6826 = ((~g3281))|((~II6825));
assign g9873 = (g9623)|(g9599)|(g9758);
assign II15759 = ((~g10267));
assign g2819 = ((~g2159));
assign g8413 = (g722&g8146);
assign g8065 = ((~II12913));
assign II12634 = ((~g7727));
assign II8677 = ((~g4374))|((~II8676));
assign II9391 = ((~g5013));
assign g6227 = ((~g5446));
assign II5539 = ((~g1270))|((~II5538));
assign g9449 = ((~g9094));
assign g6838 = (g192&g6596);
assign II10198 = ((~g6118));
assign II14330 = ((~g8819));
assign II8495 = ((~g4325));
assign II6052 = ((~g2220));
assign g3507 = ((~g3307));
assign g8526 = ((~II13735));
assign g10350 = ((~II15814));
assign g10159 = ((~II15473));
assign g5209 = ((~II8625))|((~II8626));
assign II8788 = ((~g1141))|((~II8786));
assign g2342 = ((~II5406));
assign II7131 = ((~g2640));
assign g9267 = ((~g8892));
assign g9848 = (g9724&g9557);
assign II12415 = ((~g7631));
assign g2749 = ((~II5815));
assign g6162 = (g3584&g5200);
assign g2523 = ((~II5632));
assign g8247 = (g8010)|(g7704);
assign g9925 = (g9867)|(g9712);
assign g8638 = (g8108)|(g8461);
assign II7837 = ((~g4158));
assign g10870 = ((~II16580));
assign II7899 = ((~g3380));
assign g3252 = ((~II6414));
assign II5105 = ((~g431))|((~II5104));
assign g8375 = ((~II13475));
assign g5763 = ((~g5350)&(~g5345));
assign II10237 = ((~g6120));
assign g5041 = (g3983&g4401);
assign II8085 = ((~g3664));
assign g11059 = ((~g10974));
assign II14382 = ((~g8886));
assign g8877 = (g8103&g6764&g8858);
assign g4804 = (g476&g3458);
assign g5281 = ((~g4428));
assign g2164 = ((~II5095));
assign g8301 = ((~II13266))|((~II13267));
assign g9650 = (g2797&g9240);
assign g4545 = ((~II7952));
assign g6000 = (g5480)|(g3912);
assign g2125 = ((~II5053));
assign g11485 = (g6646)|(g11462);
assign g7997 = ((~g7697));
assign g6628 = (g351&g6182);
assign g4564 = ((~g3880));
assign g5424 = ((~II8865));
assign II5414 = ((~g904));
assign g4056 = ((~II7173));
assign g10420 = ((~g10329)&(~g3744));
assign g2115 = ((~II5014))|((~II5015));
assign II15497 = ((~g10119));
assign II7984 = ((~g3621));
assign g6739 = (g5769)|(g5780);
assign g11216 = (g956&g11162);
assign II16172 = ((~g10498));
assign g4328 = ((~g4130));
assign g4606 = ((~g3829));
assign g11274 = (g4913&g11197);
assign II7938 = ((~g3406));
assign g3828 = ((~g2920));
assign II4951 = ((~g262));
assign g6112 = ((~II9789));
assign II11214 = ((~g6528));
assign II10069 = ((~g5787));
assign II6832 = ((~g2909));
assign II5204 = ((~g374))|((~II5202));
assign g10472 = ((~II16016))|((~II16017));
assign g3773 = ((~II6996));
assign g4332 = ((~g4130));
assign g9722 = (g9612)|(g9643)|(g9410)|(II14855);
assign g10378 = ((~II15858));
assign II11743 = ((~g7035));
assign II13379 = ((~g8133));
assign g7107 = ((~II11342));
assign g6099 = (g5273)|(g4550);
assign g6362 = (g5846&g4450);
assign II15362 = ((~g9987));
assign g5051 = (g4432&g2834);
assign II16209 = ((~g10452));
assign g8382 = (g6077&g8213);
assign II9531 = ((~g5004));
assign g5183 = ((~g4640));
assign g4715 = (g1077&g3638);
assign II8576 = ((~g4234))|((~II8575));
assign II15880 = ((~g2719))|((~II15878));
assign g7500 = ((~g6943));
assign g7928 = ((~g7508));
assign g6140 = ((~II9851));
assign g3757 = ((~II6952));
assign II15974 = ((~g10411));
assign II15220 = (g9841)|(g9966)|(g9857)|(g9877);
assign g9355 = ((~II14570));
assign II12060 = ((~g6961))|((~g1478));
assign g10697 = ((~II16370));
assign II5006 = ((~g421))|((~II5005));
assign g9027 = ((~II14418));
assign g5987 = ((~II9605));
assign II9984 = ((~g5529));
assign g2586 = ((~g1972));
assign g9274 = (g8974&g5708);
assign II13335 = ((~g8206));
assign II8247 = ((~g4615));
assign g7236 = (g6684)|(g6092);
assign g7295 = (g7071)|(g6321);
assign g3718 = (g192&g3164);
assign g9987 = ((~II15187));
assign g6157 = ((~II9880));
assign g6335 = ((~II10228));
assign g3804 = (g3098&g2203);
assign II7311 = ((~g2803));
assign g8702 = ((~g8664));
assign II13766 = ((~g731))|((~II13765));
assign g10547 = ((~II16206));
assign g6294 = ((~II10141));
assign g4062 = ((~II7185));
assign g6250 = ((~II10009));
assign g7795 = ((~II12550));
assign g11573 = ((~g11561));
assign g11501 = ((~II17522));
assign g10493 = ((~II16114));
assign II16376 = ((~g10596));
assign g4129 = ((~II7280));
assign g8815 = (g7948)|(g8730);
assign g11161 = (g1969&g10937);
assign g8653 = (g8526&g4013);
assign II5336 = ((~g1700));
assign II5982 = ((~g2510));
assign g8436 = ((~II13606));
assign g4116 = ((~II7260));
assign II17568 = ((~g11496))|((~II17567));
assign II10557 = ((~g6197));
assign g9707 = (g1583&g9474);
assign II7833 = ((~g3585));
assign g6050 = ((~II9677));
assign g8108 = (g1891&g7938);
assign g6745 = (g5605&g6158);
assign g7326 = ((~II11626));
assign g11268 = (g11194)|(g11030);
assign g7707 = (g691&g7206);
assign g11039 = ((~II16778));
assign II10931 = ((~g6395))|((~II10930));
assign g5151 = (g4478&g2733);
assign II15980 = ((~g10414));
assign g2943 = ((~II6125))|((~II6126));
assign g11655 = ((~II17767));
assign g9963 = (g9953&g9536);
assign g8018 = (g7742&g7425);
assign g3728 = ((~II6904));
assign g5982 = ((~II9598));
assign g4786 = ((~II8154));
assign II13595 = ((~g8339));
assign g8944 = (g8799)|(g8708);
assign g2089 = ((~II4917));
assign II5502 = ((~g1007))|((~II5500));
assign g4173 = ((~II7336));
assign g8698 = (g7591&g8576);
assign g5028 = (g4836)|(g4128);
assign II11620 = ((~g6840));
assign g9862 = (g1601&g9777);
assign g5443 = ((~II8872));
assign II8481 = ((~g3530))|((~II8479));
assign II5801 = ((~g1984));
assign II10391 = ((~g5838));
assign g7021 = ((~II11162));
assign II9077 = ((~g4765));
assign g6731 = ((~g6001));
assign II13267 = ((~g8154))|((~II13265));
assign g9584 = (g2726&g9173);
assign II13357 = ((~g8125));
assign g6406 = ((~II10314));
assign g5147 = ((~II8544))|((~II8545));
assign g9916 = (g9855)|(g9694);
assign g6298 = ((~II10153));
assign II6648 = ((~g2635));
assign g5552 = ((~g4777))|((~g4401));
assign II12574 = ((~g7522));
assign II6010 = ((~g2256));
assign II11635 = ((~g6947));
assign g8735 = (g7600&g8632);
assign II13729 = ((~g8290));
assign g3206 = ((~g2055));
assign g2744 = (II5804)|(II5805);
assign g2913 = ((~II6088));
assign II6381 = ((~g2257));
assign g8054 = (g7584&g5919);
assign g2167 = ((~II5105))|((~II5106));
assign g7535 = (g7148&g2874);
assign II16944 = ((~g11079));
assign II9099 = ((~g5572));
assign II11088 = ((~g6434));
assign II8739 = ((~g4607))|((~II8738));
assign II6867 = ((~g2949));
assign g5105 = ((~II8487));
assign g5949 = ((~II9591));
assign II12580 = ((~g7540));
assign II6531 = ((~g3186));
assign II7070 = ((~g3138));
assign g3107 = ((~g2501)&(~g2499));
assign g11600 = (g1346&g11573);
assign g4722 = (g426&g3353);
assign g4967 = (g1515&g4682);
assign II14373 = ((~g8956));
assign g5668 = ((~II9165));
assign g8281 = (g8097)|(g7818);
assign g6593 = ((~II10557));
assign g7960 = ((~g7409))|((~g5573));
assign II16111 = ((~g10385));
assign II6784 = ((~g2742));
assign II7426 = ((~g3334));
assign g2230 = ((~g704));
assign II15669 = ((~g10194));
assign II9144 = ((~g5007));
assign g11018 = (g7286&g10974);
assign g9727 = (g9650)|(g9663)|(g9362)|(II14866);
assign g6259 = ((~II10036));
assign g10160 = ((~II15476));
assign g7985 = ((~II12799));
assign II11611 = ((~g6913));
assign II16045 = ((~g833))|((~II16044));
assign II16543 = ((~g10747));
assign II17761 = ((~g11652));
assign g5288 = ((~g4438));
assign g8149 = ((~II13036));
assign g7711 = ((~II12344));
assign g6340 = ((~II10243));
assign II17052 = ((~g10923))|((~II17051));
assign g10402 = (g10295)|(g9554);
assign II11272 = ((~g6546));
assign g10269 = ((~g10154));
assign II11162 = ((~g6479));
assign g10260 = ((~g10125));
assign g8603 = (g3983&g8548);
assign g5791 = ((~II9391));
assign II6217 = ((~g2302));
assign II12790 = ((~g7618));
assign II9424 = ((~g4963));
assign g11263 = (g11187)|(g11025);
assign g8171 = ((~II13068));
assign g9364 = (g965&g9223);
assign g4608 = ((~g3829));
assign g5632 = (g1636&g4563);
assign g7586 = (g7096&g5423);
assign g4560 = (g431&g4002);
assign g3209 = ((~g2550))|((~g2061))|((~g2564))|((~g2571));
assign II4943 = ((~g324))|((~II4941));
assign g9858 = (g1595&g9774);
assign g10470 = ((~II16008))|((~II16009));
assign II17482 = ((~g11479));
assign g11631 = ((~II17707));
assign g8709 = ((~g8674));
assign g2072 = ((~II4876));
assign g9311 = ((~II14506));
assign g6902 = (g6794)|(g4223);
assign g10661 = (g10594&g3015);
assign II11204 = ((~g6523));
assign g6263 = ((~II10048));
assign g5706 = (g1574&g5121);
assign g8197 = ((~II13128));
assign II9632 = ((~g5557));
assign g8652 = (g8523&g4013);
assign II7719 = ((~g3752));
assign g7777 = ((~II12496));
assign II15452 = ((~g10058))|((~II15451));
assign II6350 = (g2445)|(g2437)|(g2433)|(g2419);
assign g10570 = ((~g10542)&(~g10324));
assign g4933 = ((~II8298));
assign g10258 = ((~g10198));
assign g8485 = ((~g8341));
assign g8647 = (g8130)|(g8470);
assign g10319 = ((~g10270));
assign g7878 = ((~g7479));
assign g2632 = ((~g2002));
assign g9536 = (g9335)|(g9331)|(g9328)|(g9324);
assign II16691 = ((~g10788));
assign g7549 = (g7269&g3829);
assign g9818 = ((~II14955));
assign g9836 = (g9737&g9785);
assign g6351 = (g6210&g5052);
assign II6535 = ((~g2826));
assign II12901 = ((~g7984));
assign g11200 = ((~g11112));
assign II11293 = ((~g6516));
assign g7442 = ((~g7237));
assign g7754 = ((~II12427));
assign g6074 = (g5349)|(g1);
assign II8805 = ((~g1113))|((~II8803));
assign g7113 = ((~II11348));
assign g5519 = ((~g4811));
assign g3862 = ((~g2920));
assign II16181 = ((~g10491));
assign g9839 = (g9702&g9742);
assign g10754 = ((~II16439));
assign g2160 = (g745&g746);
assign II13612 = ((~g8325));
assign II15461 = ((~g10074));
assign g7634 = ((~II12242));
assign g4162 = (g3106&g2971);
assign g2002 = ((~g818));
assign g8936 = (g8115&g6778&g8849);
assign g4871 = (g1864&g3523);
assign g2989 = ((~g2135));
assign g5227 = ((~II8677))|((~II8678));
assign g7848 = ((~II12641));
assign g4506 = (g1113&g3944);
assign II16008 = ((~g10424))|((~II16007));
assign g8643 = (g8364)|(g8508);
assign g10058 = ((~II15281));
assign g7883 = ((~g7689));
assign II16193 = ((~g10485));
assign g8488 = (g3664)|(g8390);
assign II10331 = ((~g6198));
assign g3393 = ((~g3144));
assign g11060 = ((~g10937));
assign g3368 = ((~g3138));
assign g10949 = (g2947&g10809);
assign g5915 = (g4168&g4977);
assign g9623 = (g17&g9274);
assign g10741 = (g10635&g4013);
assign g2602 = ((~II5707));
assign g6032 = ((~g3430)&(~g5039));
assign g2106 = ((~II4979))|((~II4980));
assign g9309 = ((~g8892));
assign II11489 = ((~g6569));
assign g2155 = ((~II5070));
assign g8141 = ((~II13020));
assign II14361 = ((~g8951));
assign g2612 = ((~II5737));
assign g9832 = ((~II14989));
assign g11462 = (g11431&g5446);
assign g11199 = ((~g11112));
assign g4549 = ((~II7956));
assign g4524 = ((~g3946));
assign g4274 = (g4054)|(g4058);
assign g5117 = ((~g4682));
assign g2244 = ((~II5251));
assign g11029 = (g401&g10974);
assign II10150 = ((~g5705));
assign II6207 = ((~g2534))|((~g802));
assign II4938 = ((~g261));
assign II12069 = ((~g139))|((~II12067));
assign g8753 = (g7414&g8664);
assign II10538 = ((~g5910));
assign g10232 = (g8892&g10150);
assign II11689 = ((~g7044));
assign g10154 = ((~II15458));
assign g5101 = ((~II8473));
assign II5528 = ((~g1265))|((~g1015));
assign II6549 = ((~g2838));
assign g3703 = ((~g2920));
assign II6137 = ((~g2496))|((~II6136));
assign II12481 = ((~g7570));
assign g9903 = (g9885&g9673);
assign g10247 = ((~II15639));
assign g5655 = ((~II9126));
assign II9317 = ((~g5576));
assign g10326 = ((~II15768));
assign g8315 = ((~II13329));
assign g8001 = ((~II12829));
assign g2653 = ((~g2011));
assign g10316 = (g10223&g9097);
assign g8959 = ((~II14326));
assign II10317 = ((~g6003));
assign g11234 = (g5424&g11106);
assign g11239 = ((~g11112));
assign g7616 = ((~II12196));
assign g8518 = ((~II13723));
assign g4478 = ((~g3820));
assign g9706 = (g9644)|(g9386)|(g9591);
assign g4989 = (g1424&g4682);
assign g6796 = ((~g6252));
assign g2956 = ((~II6159));
assign II8337 = ((~g4352));
assign g4385 = ((~II7710));
assign g8011 = ((~II12853));
assign g2418 = ((~II5497));
assign II9177 = ((~g4904));
assign g4210 = ((~II7447));
assign g6276 = ((~II10087));
assign g4372 = ((~II7677));
assign II4924 = ((~g123));
assign g3742 = ((~II6929));
assign g3538 = ((~II6726));
assign g6475 = ((~g5987));
assign g6118 = ((~II9807));
assign g6829 = (g213&g6596);
assign II5970 = ((~g2185));
assign g8121 = ((~II12978));
assign g5675 = (g131&g5361);
assign II12019 = ((~g7119))|((~g166));
assign g9611 = (g2651&g9010);
assign g5530 = (g1636&g4305);
assign g6124 = (g5181)|(g5188);
assign g6382 = ((~II10278));
assign g5774 = ((~II9362));
assign II15054 = (g7853)|(g9782)|(g9624)|(g9785);
assign g11256 = (g11186)|(g11018);
assign g4553 = (g435&g3995);
assign g2609 = ((~II5728));
assign g2774 = ((~g2276));
assign g10879 = ((~II16607));
assign g2175 = ((~g44));
assign g7244 = (g6699)|(g4720);
assign g6741 = (g3284&g6141);
assign II11519 = ((~g6591));
assign g11190 = (g5623&g11065);
assign g2881 = ((~II6031));
assign II6982 = ((~g2889));
assign g11470 = ((~II17447));
assign II16853 = ((~g10907));
assign g3633 = ((~II6802));
assign g6931 = ((~II11055));
assign g11297 = (g5490&g11242);
assign II15200 = (g9837)|(g9962)|(g9848)|(g9880);
assign g3733 = ((~II6917));
assign II6448 = ((~g2264))|((~II6447));
assign g4428 = ((~II7776));
assign g2758 = ((~II5840));
assign g9223 = (g6454&g8960);
assign g10505 = ((~g10432))|((~g5938));
assign II6391 = ((~g2478));
assign II14979 = ((~g9671));
assign g2645 = ((~g1991));
assign g10760 = (g10695&g10691);
assign II6347 = ((~g2462));
assign II12115 = ((~g162))|((~II12113));
assign g10737 = (g10687&g4840);
assign g5012 = ((~II8388));
assign II17764 = ((~g11651));
assign g2124 = ((~II5050));
assign g3876 = ((~II7061));
assign g7745 = ((~II12400));
assign g8563 = ((~II13782));
assign g5256 = (g4297&g2779);
assign II5421 = ((~g549));
assign g8133 = ((~II13002));
assign II16670 = ((~g10797));
assign II16108 = ((~g10383));
assign g8806 = (g7931)|(g8718);
assign II12205 = ((~g6993));
assign g10792 = ((~II16492));
assign g9874 = ((~g9519)&(~g9536)&(~g9579)&(~II15033));
assign g3735 = ((~II6921));
assign g2971 = ((~g2046));
assign g8720 = (g8601&g7905);
assign g6199 = (g557&g5062);
assign II8614 = ((~g4414));
assign II6183 = ((~g2131));
assign II13545 = ((~g713))|((~II13544));
assign g6704 = ((~g5949));
assign g4914 = (g1062&g4436);
assign II13457 = ((~g8184));
assign II6240 = ((~g878));
assign II17365 = ((~g11380));
assign II7760 = ((~g3768));
assign II6188 = ((~g466))|((~II6186));
assign g6133 = ((~II9836));
assign II12046 = ((~g6951))|((~II12045));
assign II5240 = ((~g64));
assign g8400 = (g6097&g8234);
assign g9489 = ((~g9052)&(~g9030));
assign g11194 = (g5637&g11067);
assign II8865 = ((~g4518));
assign II15215 = (g9840)|(g9965)|(g9854)|(g9879);
assign II6247 = ((~g2462));
assign g4681 = ((~g3546));
assign g6439 = (g4479&g5919);
assign g9345 = ((~II14540));
assign g6213 = ((~g5426));
assign g11326 = (g11296)|(g11166);
assign g8024 = (g7394&g4337);
assign g9846 = (g287&g9764);
assign g4819 = ((~g3354));
assign g3142 = ((~II6360));
assign II6398 = ((~g2335));
assign g2826 = ((~g2163));
assign II7680 = ((~g3736));
assign II7064 = ((~g2984));
assign g6844 = ((~II10904));
assign g6893 = ((~II10991));
assign g11290 = (g11246&g4226);
assign g10857 = (g6090)|(g10738);
assign g9572 = ((~II14709));
assign II7244 = ((~g3226));
assign g11411 = ((~II17274));
assign II14080 = ((~g8714));
assign II15491 = ((~g10093));
assign g5745 = (g1549&g5192);
assign II5031 = ((~g928));
assign II13791 = ((~g8518));
assign II14265 = ((~g1814))|((~II14263));
assign g11105 = (g3634&g10937);
assign g3513 = (g3118)|(g2180);
assign g7305 = ((~II11563));
assign g11414 = ((~II17282))|((~II17283));
assign g2939 = (g2411&g1687);
assign g8967 = (g8085&g6778&g8849);
assign g7512 = ((~g7148));
assign g8631 = (g8474)|(g7449);
assign II17687 = ((~g11610));
assign g6057 = ((~g5446));
assign g6571 = ((~II10503));
assign g2208 = ((~g84));
assign g6447 = ((~g6166));
assign g8511 = ((~g5277))|((~g8366));
assign II11043 = ((~g6412));
assign g2045 = ((~g1811));
assign g7110 = ((~II11345));
assign g5637 = ((~II9074));
assign g1969 = ((~g456));
assign g2916 = ((~II6097));
assign g3751 = ((~II6944));
assign g10501 = (g4161)|(g10445);
assign II7556 = ((~g4080));
assign II5952 = ((~g2506));
assign II5450 = ((~g1235))|((~II5449));
assign g4471 = (g1121&g3862);
assign g10115 = ((~II15353));
assign g2446 = ((~g1400));
assign g10937 = (g4822&g10822);
assign g7947 = ((~g7395))|((~g7390))|((~g7279))|((~g7369));
assign II15672 = ((~g10132));
assign g8310 = ((~II13314));
assign g7453 = (g7148&g2809);
assign g8795 = ((~II14112));
assign g8960 = (g8085&g6368&g8828);
assign g10720 = (g10304)|(g10667);
assign g8338 = ((~II13394));
assign g5880 = ((~g5361));
assign g10863 = (g5531)|(g10750);
assign g3905 = ((~g2920));
assign II7973 = ((~g3437));
assign g8333 = ((~II13379));
assign II12354 = ((~g7143));
assign g9927 = (g9869)|(g9716);
assign g8623 = ((~II13877))|((~II13878));
assign g5308 = ((~II8787))|((~II8788));
assign g8276 = ((~II13200));
assign g8295 = ((~II13239));
assign g6824 = (g1371&g6596);
assign g4353 = ((~II7636));
assign II6944 = ((~g2859));
assign g2544 = (g1341&g1336);
assign g6870 = ((~II10952));
assign II7752 = ((~g3407));
assign II4996 = ((~g416))|((~II4995));
assign g11067 = ((~g10974));
assign II6560 = ((~g2845));
assign II6323 = ((~g2050))|((~II6322));
assign II17752 = ((~g11645));
assign g11599 = (g1341&g11572);
assign II5676 = ((~g1218))|((~II5675));
assign II16060 = ((~g10372))|((~II16058));
assign g9920 = (g9860)|(g9701);
assign II5830 = ((~g2067));
assign II11143 = ((~g6446));
assign II6924 = ((~g2843));
assign g10897 = ((~g10827));
assign II14976 = ((~g9670));
assign II12268 = ((~g7107));
assign g4511 = ((~g3586));
assign II5352 = (g1129)|(g1125)|(g1121)|(g1117);
assign g7431 = ((~II11821));
assign II6715 = ((~g2961))|((~II6714));
assign g7315 = ((~II11593));
assign g7285 = ((~II11531));
assign II15470 = ((~g10111));
assign g5112 = ((~g4682));
assign g7497 = ((~g7148));
assign g7683 = ((~g7148));
assign g3971 = ((~II7104));
assign g5813 = (g5617)|(g4869);
assign g10525 = ((~g10499));
assign g11048 = ((~II16805));
assign g10930 = ((~g10827));
assign g8924 = ((~II14249));
assign g4265 = ((~g3664));
assign g7732 = (g6935&g3880);
assign II10051 = ((~g5702));
assign g2008 = ((~g971));
assign g4920 = ((~II8293));
assign g5670 = ((~II9171));
assign g7957 = (g2885&g7527);
assign g3055 = ((~g2135));
assign g5594 = ((~II9016));
assign g4287 = ((~II7546));
assign II13554 = ((~g8262))|((~II13552));
assign II6818 = ((~g2758));
assign II16031 = ((~g829))|((~II16030));
assign g10769 = (g10652&g4840);
assign II14675 = ((~g9263));
assign g7916 = ((~g7651));
assign g2563 = (II5689&II5690);
assign g6172 = ((~II9901));
assign g11604 = (g11583)|(g11554);
assign II6572 = ((~g2853));
assign g11286 = (g10670)|(g11209);
assign g5603 = ((~II9029));
assign g7140 = (g6069&g6711);
assign g4399 = ((~g3638));
assign II5317 = ((~g1027))|((~II5315));
assign g6621 = (g52&g6164);
assign II16016 = ((~g10425))|((~II16015));
assign g5738 = (g1586&g5184);
assign g10356 = ((~II15832));
assign g2834 = ((~II5952));
assign g8260 = (g2775&g7911);
assign g7344 = ((~II11680));
assign g11094 = (g374&g10883);
assign g6243 = (g5537)|(g4774);
assign II7600 = ((~g4159));
assign g9450 = ((~g9097));
assign g11366 = ((~II17191));
assign g6468 = (g5690)|(g4950);
assign g7141 = (g6073&g6716);
assign g11030 = (g406&g10974);
assign g3473 = ((~II6676));
assign g11087 = (g829&g10950);
assign g2067 = ((~g108));
assign g2196 = ((~g91));
assign II7697 = ((~g3743));
assign g10970 = (g10852&g3390);
assign II13773 = ((~g8384));
assign g2012 = ((~g981));
assign g6673 = (g5305&g5822);
assign g10646 = (g10625)|(g7739);
assign g8233 = ((~g7872));
assign II11961 = ((~g7053));
assign g7362 = ((~II11734));
assign II14933 = ((~g9454));
assign g2845 = ((~g2168));
assign g7145 = (g6082&g6718);
assign II14176 = ((~g8784));
assign g11008 = (g5171&g10827);
assign g11346 = ((~II17161));
assign II16311 = ((~g10584));
assign g10702 = (g10562)|(g3877);
assign II14405 = ((~g8937));
assign g9948 = (g9928&g9392);
assign g7661 = (g7127&g2251);
assign g2751 = ((~II5821));
assign g8930 = (g8100&g6368&g8828);
assign g4895 = ((~II8250));
assign g11543 = ((~g11519));
assign g7047 = ((~II11222));
assign g6886 = (g1932&g6420);
assign g4941 = (g1038&g4451);
assign II14534 = ((~g9290));
assign g7877 = ((~g7479));
assign g6084 = ((~II9731));
assign g10272 = ((~g10168));
assign II10009 = ((~g5542));
assign II12568 = ((~g7502));
assign g10896 = ((~II16650));
assign II6779 = ((~g650))|((~II6777));
assign II9362 = ((~g5013));
assign II5827 = ((~g2271));
assign g11611 = ((~II17657));
assign g10386 = ((~II15879))|((~II15880));
assign g10167 = ((~II15497));
assign II5929 = ((~g2225));
assign g2272 = ((~II5316))|((~II5317));
assign II16682 = ((~g10799));
assign II16796 = ((~g11016));
assign II7034 = ((~g3089))|((~II7033));
assign g6345 = (g5823&g4426);
assign II15530 = ((~g10107));
assign g2229 = ((~g162));
assign II15258 = ((~g9980))|((~II15256));
assign g5695 = (g166&g5361);
assign II10514 = ((~g6154));
assign II9065 = ((~g4760));
assign g7648 = ((~II12255));
assign II8877 = ((~g4421));
assign II11412 = ((~g6411));
assign g8282 = (g8101)|(g7819);
assign g5260 = (g1092&g4758);
assign II5995 = ((~g2196));
assign g3623 = ((~II6761))|((~II6762));
assign g6329 = (g1265&g5949);
assign g5628 = ((~II9062));
assign g7139 = (g6060&g6709);
assign g4501 = ((~g3946));
assign g7940 = (g7620&g4013);
assign g10592 = ((~II16261));
assign II17525 = ((~g11486));
assign g10330 = ((~II15778));
assign g6859 = ((~II10937));
assign g6287 = ((~II10120));
assign g10776 = (g5544)|(g10758);
assign g3496 = ((~II6686));
assign g2405 = ((~II5485))|((~II5486));
assign g7598 = ((~II12137))|((~II12138));
assign g5822 = ((~g5320));
assign II6962 = ((~g2791));
assign g11171 = (g481&g11112);
assign II9237 = ((~g5205));
assign g11403 = ((~II17252));
assign g7591 = ((~II12103));
assign g10455 = ((~II15956));
assign g9259 = ((~g8892));
assign g6863 = ((~g6740));
assign II17124 = ((~g11232));
assign II5297 = ((~g798))|((~II5295));
assign II16286 = ((~g10540));
assign g9660 = (g1188&g9125);
assign g11453 = ((~II17416));
assign g6521 = ((~II10437));
assign g7809 = ((~II12592));
assign II15907 = ((~g6899))|((~II15906));
assign II15691 = ((~g10233));
assign g9765 = ((~II14910));
assign g3040 = ((~g2135));
assign II9165 = ((~g5037));
assign g4584 = (g3710&g2322);
assign g11262 = (g11240)|(g11024);
assign g3540 = ((~g3307));
assign II13344 = ((~g8121));
assign g4065 = ((~g2794));
assign II14272 = ((~g1822))|((~II14270));
assign g4239 = (g4000)|(g4008);
assign II12846 = ((~g7685));
assign g5757 = (g1552&g5203);
assign g5350 = ((~g4163)&(~g4872));
assign g5475 = ((~II8892));
assign g10827 = ((~II16543));
assign g8041 = (g7524&g5128);
assign II10693 = ((~g6068));
assign g3769 = ((~II6982));
assign g10626 = (g10547&g4558);
assign g7079 = ((~II11312));
assign II12939 = ((~g7977));
assign g4630 = ((~g3077)&(~g3491)&(~g3485)&(~g3479));
assign g3007 = ((~II6240));
assign g5545 = (g1730&g4321);
assign g10746 = (g10643&g4013);
assign g5199 = (g1068&g4719);
assign g6623 = (g55&g6170);
assign g6184 = ((~II9915));
assign g5780 = ((~g2112)&(~g4921));
assign g8765 = (g8630&g5151);
assign II7330 = ((~g3761));
assign g8356 = ((~II13448));
assign II11262 = ((~g6775))|((~II11261));
assign g8559 = (g8380)|(g4731);
assign g4365 = ((~g3880));
assign II17416 = ((~g11420));
assign II11644 = ((~g6970));
assign g6681 = ((~g5830));
assign g5568 = ((~II8985));
assign II15347 = ((~g9995));
assign g4228 = ((~g3914));
assign g6776 = (g5809&g4390);
assign g4491 = ((~g3546));
assign II14831 = (g9613)|(g9622)|(g9586);
assign g3913 = ((~g2920));
assign g5279 = (g1766&g4783);
assign II15482 = ((~g10115));
assign g8296 = ((~II13242));
assign g6179 = (g5115&g5354);
assign g7522 = ((~II11904));
assign g8542 = ((~g2571))|((~g1828))|((~g1814))|((~g8390));
assign II12126 = ((~g7103))|((~g170));
assign II9617 = ((~g5405));
assign g6692 = ((~II10659));
assign II12153 = ((~g6874));
assign g9690 = (g266&g9432);
assign II15039 = (g7853)|(g9809)|(g9624)|(g9785);
assign g8444 = ((~II13630));
assign g9579 = (g9052)|(g9030);
assign g5219 = ((~II8651))|((~II8652));
assign g6056 = ((~g5426));
assign g5344 = ((~II8811));
assign g3715 = ((~g2920));
assign g6687 = (g5486&g5840);
assign g10900 = ((~II16656));
assign g11072 = ((~g10913));
assign g10907 = ((~II16673));
assign g10363 = ((~g10355)&(~g3566));
assign g9387 = ((~g9010)&(~g9240)&(~g9223)&(~II14596));
assign g9669 = ((~g9392)&(~g9367));
assign II13521 = ((~g695))|((~g8249));
assign g8074 = (g718&g7826);
assign g4757 = ((~II8109));
assign g7769 = ((~II12472));
assign g2017 = ((~g1218));
assign II12186 = ((~g7264));
assign g10808 = (g10744&g3829);
assign g3321 = ((~II6484));
assign g10079 = ((~II15305));
assign g4418 = ((~II7760));
assign II11879 = ((~g6893));
assign g2132 = (g1872&g1882);
assign g11333 = (g11274)|(g11173);
assign g9342 = ((~II14531));
assign II10966 = ((~g6561));
assign II5013 = ((~g1007))|((~g1011));
assign g4354 = ((~II7639));
assign II6469 = ((~g2479))|((~II6467));
assign g9652 = (g953&g9223);
assign g9269 = (g8933&g3413);
assign g7930 = (g7621&g3110);
assign II14397 = ((~g8888));
assign g7101 = ((~g6617))|((~g2364));
assign g10558 = (g4126)|(g10510);
assign II9040 = ((~g4794));
assign II15476 = ((~g10114));
assign g5521 = ((~g4530));
assign g7038 = ((~II11201));
assign g8983 = ((~II14370));
assign II6330 = (g2549&g2556&g2562&g2570);
assign g10597 = (g10533&g4359);
assign g11518 = ((~II17563));
assign II10920 = ((~g6733));
assign g4379 = ((~g3698));
assign II12380 = ((~g7204));
assign g3622 = ((~II6757));
assign II16264 = ((~g10557));
assign II17400 = ((~g11418))|((~g11416));
assign II16088 = ((~g10375))|((~II16086));
assign g4617 = (g3275&g3879);
assign g5734 = ((~II9290));
assign II13013 = ((~g8048));
assign II10030 = ((~g5685));
assign g7939 = (g2829&g7460);
assign g6533 = (g5771)|(g5002);
assign g6190 = ((~g5426));
assign g4123 = (g2695&g3037);
assign g11100 = (g853&g10950);
assign g10136 = ((~II15406));
assign g4724 = ((~g3586));
assign II14822 = (g9597)|(g9604)|(g9582);
assign g9934 = (g9913&g9624);
assign g2525 = (g762&g758);
assign g3407 = (g2561&g3012);
assign g2242 = ((~II5245));
assign g5993 = (g5090)|(g4400);
assign II15072 = ((~g9713));
assign g5824 = (g5602)|(g4839);
assign g8225 = ((~g7826));
assign g5262 = ((~g4353));
assign g4187 = ((~II7378));
assign g3334 = ((~II6517));
assign g6657 = ((~II10620));
assign II7002 = ((~g2907));
assign II8889 = ((~g4553));
assign g5422 = ((~g4470));
assign II13403 = ((~g8236));
assign g7351 = ((~II11701));
assign g11594 = ((~II17636));
assign g8102 = (g6209&g7878);
assign II7923 = ((~g3394));
assign g9741 = ((~II14888));
assign g8313 = ((~II13323));
assign g5744 = (g1528&g5191);
assign g11513 = ((~II17558));
assign g6645 = (g67&g6202);
assign g3628 = ((~g3111));
assign g6984 = ((~g6382));
assign g5576 = (g4675)|(g3664);
assign II5913 = ((~g2169));
assign g8448 = ((~II13642));
assign g8364 = (g658&g8235);
assign g2060 = ((~g1380));
assign g6023 = ((~g2763)&(~g4975));
assign II6019 = ((~g2554));
assign II12592 = ((~g7445));
assign g4001 = ((~g3200));
assign g9264 = ((~II14477));
assign g8722 = (g8604&g7908);
assign g6400 = ((~II10308));
assign g4305 = ((~g4013));
assign g9821 = ((~II14964));
assign g9883 = ((~II15060));
assign II11995 = ((~g7107))|((~g127));
assign g7430 = ((~g7221));
assign g6316 = (g1270&g5949);
assign g9608 = (g7&g9292);
assign g7211 = (g6647)|(g6067);
assign g6635 = ((~II10592));
assign II10888 = ((~g6333));
assign II10520 = ((~g6231))|((~II10519));
assign g6957 = ((~II11109));
assign g10562 = ((~g10483)&(~g10529));
assign II17240 = ((~g11395));
assign g7044 = ((~II11217));
assign g6555 = ((~g5740));
assign g2753 = ((~II5827));
assign II13233 = ((~g8265));
assign II7414 = ((~g4156));
assign g10104 = ((~II15338));
assign g4838 = (g3275&g4122);
assign g7671 = ((~g7011))|((~g6995))|((~g6984))|((~g6974));
assign II15900 = ((~g10287))|((~II15898));
assign g7949 = ((~g7422));
assign g6926 = ((~II11046));
assign II13301 = ((~g1936))|((~II13300));
assign g7097 = ((~II11330));
assign g6280 = ((~II10099));
assign g5698 = (g1571&g5116);
assign g4420 = ((~II7766));
assign g3533 = (g1981&g2892);
assign g10173 = ((~g10120));
assign g6877 = ((~II10963));
assign II17419 = ((~g11421));
assign g6480 = (g5721)|(g4971);
assign II10024 = ((~g5700));
assign g10039 = ((~II15244));
assign g2852 = ((~II5982));
assign g8742 = (g8135)|(g8598);
assign II10117 = ((~g6241));
assign II4972 = ((~g991))|((~II4971));
assign g7601 = ((~II12153));
assign II6772 = ((~g382))|((~II6770));
assign g11351 = ((~II17170));
assign g9714 = (g9664)|(g9366)|(g9654);
assign g9331 = (g8972&g5708);
assign g4543 = ((~g3946));
assign II11306 = ((~g6731));
assign g10375 = ((~g10288)&(~g3463));
assign II13421 = ((~g8200));
assign II14645 = ((~g9088));
assign g2824 = ((~II5932));
assign g3287 = (g802&g2534);
assign g7065 = ((~II11272));
assign II13131 = ((~g7979));
assign II13478 = ((~g8191));
assign g3433 = ((~II6648));
assign II14776 = (g8995)|(g9205)|(g9192);
assign II15467 = ((~g10079));
assign II9159 = ((~g5033));
assign g10192 = ((~II15554));
assign g4393 = ((~II7726));
assign g9726 = (g9411)|(g9420)|(g9489);
assign g8325 = ((~II13357));
assign g7983 = ((~II12793));
assign II9007 = ((~g4492))|((~II9006));
assign g10369 = (g10361&g3382);
assign II13351 = ((~g8214));
assign II11602 = ((~g6833));
assign II15510 = ((~g10035));
assign g5417 = ((~II8854));
assign II17231 = ((~g11303));
assign g9508 = ((~g9271));
assign g4760 = (g486&g3393);
assign g7625 = (g673&g7085);
assign II7906 = ((~g3907));
assign II6938 = ((~g2854));
assign II12145 = ((~g158))|((~II12143));
assign II6806 = ((~g3268))|((~II6805));
assign g6567 = ((~II10495));
assign g8097 = (g6200&g7851);
assign g10887 = ((~II16623));
assign II12242 = ((~g7089));
assign g7779 = ((~II12502));
assign g10480 = ((~II16066))|((~II16067));
assign II11929 = ((~g6901));
assign g3365 = ((~II6553));
assign II8265 = ((~g4602));
assign II15890 = ((~g853))|((~g10286));
assign II7931 = ((~g3624));
assign g2578 = ((~g1962));
assign II6176 = ((~g2177))|((~g197));
assign II11201 = ((~g6522));
assign g7988 = (g1878&g7379);
assign g6076 = ((~II9717));
assign g11559 = (g2719&g11519);
assign g4959 = (g1520&g4682);
assign II10108 = ((~g5743));
assign g11213 = (g947&g11157);
assign II13294 = ((~g1882))|((~II13293));
assign g4341 = (g339&g3586);
assign g9945 = (g9925&g9392);
assign g8549 = ((~g5527))|((~g8390));
assign II5909 = ((~g2207));
assign g9867 = (g1552&g9807);
assign g11246 = (g11094)|(g10948);
assign g5497 = (g4296&g3522);
assign g3274 = ((~II6454));
assign II5604 = ((~g1149))|((~g1153));
assign g8303 = ((~g8209)&(~g4811));
assign g9888 = (g9648)|(g9608)|(g9757);
assign II7630 = ((~g3524));
assign II5363 = (g1149)|(g1153)|(g1157)|(g1160);
assign g7221 = ((~II11459));
assign g7802 = ((~II12571));
assign g2812 = ((~g2158));
assign g5768 = ((~II9352));
assign g6562 = ((~g5774));
assign g7743 = (g6967&g3880);
assign II13397 = ((~g8138));
assign g5684 = ((~II9205));
assign g5067 = (g305&g4811);
assign g3267 = ((~II6439));
assign g2220 = ((~g104));
assign II10770 = ((~g5944))|((~II10769));
assign II12779 = ((~g7608));
assign g7313 = ((~II11587));
assign g8430 = (g8386)|(g8070);
assign II14133 = ((~g8772));
assign g4310 = ((~II7577));
assign g6550 = (g1231&g6089);
assign II11882 = ((~g6895));
assign II13583 = ((~g8344));
assign g8158 = (g7893)|(g6883);
assign g5856 = ((~g5245));
assign g8067 = ((~II12919));
assign g8241 = (g7536)|(g7989);
assign g8575 = ((~II13816));
assign II5725 = ((~g2079));
assign II14210 = ((~g8824))|((~II14209));
assign g8478 = ((~II13678));
assign g6215 = (g1504&g5128);
assign g10296 = ((~II15708));
assign II12694 = ((~g7374));
assign II13076 = ((~g1872))|((~g7963));
assign g6499 = ((~g5867));
assign g7567 = ((~II12020))|((~II12021));
assign II10671 = ((~g6045));
assign II11629 = ((~g6914));
assign g2090 = ((~II4920));
assign g11202 = ((~g11112));
assign g11391 = (g11275&g7912);
assign II8815 = ((~g4471));
assign g3682 = ((~g2920));
assign g8443 = ((~II13627));
assign g5223 = ((~g4640));
assign g4334 = (g1160&g3703);
assign g6619 = (g49&g6156);
assign g3422 = (g225&g3228);
assign g3272 = ((~g2450));
assign g9107 = ((~II14443))|((~II14444));
assign g8595 = ((~II13840));
assign II16086 = ((~g861))|((~g10375));
assign g8875 = (g8255&g6368&g8858);
assign g2516 = ((~II5612))|((~II5613));
assign g6914 = ((~II11024));
assign II14421 = ((~g8944));
assign II5565 = ((~g1713));
assign g8798 = ((~II14119));
assign II17516 = ((~g11483));
assign II12093 = ((~g6944))|((~II12092));
assign II13091 = ((~g1840))|((~II13089));
assign II10566 = ((~g5904));
assign g2569 = ((~II5695));
assign g8348 = ((~II13424));
assign g11338 = (g11283)|(g11178);
assign g3523 = ((~g2971));
assign II15157 = ((~g9931));
assign II15616 = ((~g10043))|((~II15615));
assign g7119 = ((~II11354));
assign II17672 = ((~g11605));
assign g10262 = ((~g10142));
assign g7547 = ((~II11974))|((~II11975));
assign g5704 = (g143&g5361);
assign g11436 = ((~II17359));
assign II5251 = ((~g1424));
assign g10468 = ((~II16000))|((~II16001));
assign g7632 = (g7184&g5574);
assign II17494 = ((~g3623))|((~II17492));
assign g3970 = (g225&g3164);
assign g11182 = ((~II16947));
assign g6910 = (g6341)|(g5680);
assign g8778 = (g8688&g2317);
assign g3771 = ((~II6989))|((~II6990));
assign g6809 = ((~II10837));
assign g2117 = ((~II5024))|((~II5025));
assign g4058 = (g2707&g2276);
assign g6716 = ((~g5949));
assign g3391 = ((~g2896));
assign g2420 = ((~g237));
assign II6403 = ((~g2337));
assign II8811 = ((~g4465));
assign II16101 = ((~g10381));
assign g8820 = (g8705&g5422);
assign g8784 = ((~II14087));
assign g4550 = (g342&g3586);
assign g8529 = ((~II13738));
assign II17486 = ((~g11384))|((~II17485));
assign g10785 = (g10728&g5177);
assign g7402 = ((~g6860));
assign g7425 = ((~g7214));
assign g4537 = (g444&g3988);
assign g11442 = ((~II17377));
assign II11953 = ((~g6907));
assign g11272 = (g5629&g11193);
assign g10725 = (g4962)|(g10634);
assign g2803 = ((~g2154));
assign g5849 = (g4949)|(g4260);
assign g7082 = ((~II11315));
assign g5653 = ((~II9120));
assign g8803 = ((~II14130));
assign g4453 = ((~II7810));
assign II14967 = ((~g9763));
assign g5287 = (g3876&g4782);
assign g22 = ((~II4777));
assign II7612 = ((~g3817));
assign g8275 = ((~II13197));
assign g10583 = (g10518&g10515);
assign g11487 = (g6662)|(g11464);
assign II9446 = ((~g5052));
assign II17155 = ((~g11310));
assign II15639 = ((~g10179));
assign II15609 = ((~g10144))|((~II15607));
assign II5424 = ((~g910));
assign g4515 = ((~II7916));
assign II4876 = ((~g580));
assign g2790 = ((~g2276));
assign II6881 = ((~g1351))|((~II6879));
assign g6126 = (g5639&g4319);
assign g8249 = (g8018)|(g7710);
assign II9734 = ((~g5257));
assign g4802 = ((~g3337));
assign g4258 = ((~II7509));
assign g11254 = (g986&g11073);
assign g3662 = ((~II6826))|((~II6827));
assign g9774 = ((~g9474));
assign II9826 = ((~g5390));
assign g6451 = ((~II10381));
assign g8712 = ((~g8680));
assign g11057 = ((~g10937));
assign II15199 = (g8167)|(g9903)|(g9932)|(g9828);
assign g11287 = ((~g11207));
assign g7054 = ((~II11242))|((~II11243));
assign g10145 = ((~II15437));
assign g8758 = ((~II14055));
assign II8786 = ((~g4639))|((~g1141));
assign g2267 = ((~II5304));
assign g8477 = ((~g8317));
assign II15795 = ((~g10280));
assign II9216 = ((~g4935));
assign g4970 = ((~g4411));
assign g3093 = ((~II6299));
assign II7864 = ((~g4099))|((~II7863));
assign g4489 = (g348&g3586);
assign g8046 = (g7548&g5128);
assign g5618 = (g1630&g4551);
assign g2539 = ((~II5652));
assign g7826 = ((~II12627));
assign g3505 = ((~II6694));
assign g11464 = (g11433&g5446);
assign g4639 = ((~g3501)&(~g2669)&(~g2662)&(~g2655));
assign g4326 = ((~g3863));
assign g5390 = (g3220&g4819);
assign g8671 = ((~II13956));
assign g10183 = ((~g10042));
assign II14326 = ((~g8818));
assign g2713 = ((~g2042));
assign II15079 = ((~g9745));
assign g9429 = ((~g9082));
assign g2085 = ((~II4903));
assign g2962 = ((~II6183));
assign g8613 = ((~g8484));
assign II7840 = ((~g3431));
assign g10473 = ((~g10380));
assign II15507 = ((~g10047));
assign g10394 = ((~II15899))|((~II15900));
assign g3138 = ((~II6356));
assign g7395 = ((~g6941));
assign II14355 = ((~g8948));
assign II5858 = ((~g2529));
assign g9842 = (g9708&g9516);
assign g6708 = ((~II10689));
assign g5200 = ((~g4567));
assign II8089 = ((~g3545));
assign II9564 = ((~g5109));
assign II12214 = ((~g7061))|((~g2518));
assign II16546 = ((~g10724));
assign g10715 = (g2272&g10630);
assign II16574 = ((~g10821));
assign II5530 = ((~g1015))|((~II5528));
assign II6199 = ((~g2525))|((~g766));
assign II12138 = ((~g131))|((~II12136));
assign II12445 = ((~g7521));
assign II12867 = ((~g7638));
assign g5084 = (g1776&g4591);
assign II17289 = ((~g11366))|((~II17288));
assign II16589 = ((~g10820));
assign II10325 = ((~g6003));
assign II9329 = ((~g5504));
assign g4480 = (g1133&g3905);
assign II6654 = ((~g2952));
assign g9676 = (g9454)|(g9292)|(g9274);
assign g3328 = ((~II6501));
assign g6513 = (g5737)|(g4991);
assign g7750 = ((~II12415));
assign II12171 = ((~g6885));
assign II12451 = ((~g7538));
assign g4572 = ((~g3419)&(~g3408)&(~g3628));
assign II10531 = ((~g6169));
assign g2345 = ((~g1936));
assign g7999 = ((~II12825));
assign g8343 = ((~II13409));
assign g9893 = ((~II15082));
assign g4784 = (g506&g3432);
assign g10253 = ((~g10138));
assign II9695 = ((~g5212));
assign g7904 = ((~II12690));
assign II11280 = ((~g6485))|((~II11278));
assign II6428 = ((~g2348));
assign g9871 = (g1564&g9668);
assign g11644 = ((~II17736));
assign II16187 = ((~g10492));
assign II13514 = ((~g686))|((~II13513));
assign g5232 = ((~g4640));
assign II11889 = ((~g6898));
assign II5044 = ((~g1182));
assign g10498 = ((~II16121));
assign g6938 = ((~II11068));
assign II9731 = ((~g5255));
assign g5192 = ((~g4640));
assign II11333 = ((~g6670));
assign g6789 = ((~II10789));
assign II8551 = ((~g4342));
assign II5047 = ((~g1185));
assign II12289 = ((~g7142));
assign g8176 = (g5299&g7853);
assign g8738 = ((~g8688))|((~g4921));
assign II7348 = ((~g4056));
assign g11657 = ((~II17773));
assign g5641 = ((~II9084));
assign g10481 = ((~II16073))|((~II16074));
assign g10469 = ((~g10430))|((~g5999));
assign II11222 = ((~g6533));
assign II9229 = ((~g4954));
assign II16580 = ((~g10826));
assign g5840 = ((~g5320));
assign g7724 = ((~II12357));
assign g10451 = (g10444&g3365);
assign II13978 = ((~g8575));
assign g10619 = ((~II16292));
assign g4567 = ((~g3374));
assign g9670 = ((~II14799));
assign g11629 = ((~II17701));
assign II11821 = ((~g7205));
assign II16307 = ((~g10589));
assign g7816 = ((~II12613));
assign g10752 = (g10692&g3586);
assign g7329 = ((~II11635));
assign g6241 = ((~II9992));
assign g8755 = (g7426&g8671);
assign g5127 = ((~II8535));
assign g2437 = ((~II5529))|((~II5530));
assign g11186 = (g5594&g11059);
assign g1980 = ((~g646));
assign g2742 = ((~II5798));
assign g5837 = (g5640)|(g4224);
assign g2165 = ((~II5098));
assign g6752 = (g6187&g2343);
assign g8570 = ((~II13803));
assign g2988 = ((~II6225))|((~II6226));
assign II13326 = ((~g8203));
assign g4881 = (g991&g3914);
assign g10522 = ((~g10486)&(~g10239));
assign II6043 = ((~g2267));
assign II7216 = ((~g2952));
assign II11242 = ((~g6760))|((~II11241));
assign g8605 = (g8404)|(g8553);
assign II9574 = ((~g5608))|((~g818));
assign II5067 = ((~g33));
assign II8259 = ((~g4590));
assign g11406 = ((~II17261));
assign g10239 = ((~g9317)&(~g10179));
assign g11446 = ((~II17387));
assign g5528 = (g4322&g3537);
assign g5078 = ((~g4372));
assign g11425 = (g11350&g10899);
assign g8185 = (g664&g7997);
assign II5165 = ((~g1508))|((~II5164));
assign II12397 = ((~g7284));
assign g3982 = ((~g3052));
assign II7009 = ((~g2913));
assign II9842 = ((~g5405));
assign g2099 = ((~II4942))|((~II4943));
assign g2994 = ((~g2057));
assign g8719 = ((~g8579));
assign g5397 = ((~II8835));
assign II8147 = ((~g3633));
assign g3816 = ((~g3228));
assign g11015 = (g5217&g10827);
assign II11459 = ((~g6488));
assign II6097 = ((~g2391));
assign II10286 = ((~g6237));
assign g6797 = ((~II10801));
assign g7051 = ((~II11232));
assign g2391 = ((~II5478));
assign g10206 = ((~g10178));
assign g8161 = (g8005)|(g7185);
assign II7886 = ((~g4076));
assign g4466 = ((~II7833));
assign g4295 = ((~II7556));
assign g5172 = (g4555&g4549);
assign II5089 = ((~g1854));
assign g2562 = ((~g1383));
assign II6702 = ((~g2801));
assign g7785 = ((~II12520));
assign g6238 = (g572&g5096);
assign g8629 = ((~II13901))|((~II13902));
assign g3260 = ((~II6428));
assign g6790 = (g5813&g4398);
assign g4204 = ((~II7429));
assign II11509 = ((~g6580))|((~II11508));
assign g3359 = ((~II6543));
assign g3104 = (II6316&II6317);
assign g7685 = ((~g7148));
assign g97 = ((~II4780));
assign g2797 = ((~g2524));
assign g7783 = ((~II12514));
assign g5912 = ((~II9544));
assign g4737 = ((~g3440));
assign g7389 = (g7001&g3880);
assign II11967 = ((~g6911));
assign II10352 = ((~g6216));
assign II14127 = ((~g8768));
assign II13265 = ((~g1909))|((~g8154));
assign g4816 = (g4070&g2336);
assign g6713 = ((~II10698));
assign g5360 = ((~g2071)&(~g4225));
assign g2206 = ((~II5171));
assign g7686 = ((~g7148));
assign g6807 = ((~II10831));
assign g7955 = (g2877&g7516);
assign II16781 = ((~g10893));
assign g2198 = ((~g668));
assign g10712 = (g10662)|(g9531);
assign II15811 = ((~g10200));
assign g5672 = ((~II9177));
assign II16739 = ((~g10856));
assign g9348 = ((~II14549));
assign II7858 = ((~g3631));
assign g11409 = ((~II17268));
assign g9647 = ((~g9125)&(~g9111)&(~g9173)&(~g9151));
assign g10533 = (g4933)|(g10449);
assign g8350 = ((~II13430));
assign g5605 = (g4828&g704);
assign g8289 = (g6777&g8109&g6475);
assign II7096 = ((~g3186));
assign g8659 = (g8535&g4013);
assign II9863 = ((~g5557));
assign g6646 = (g360&g6203);
assign g10110 = ((~II15344));
assign II6807 = ((~g471))|((~II6805));
assign II12604 = ((~g7630));
assign g2479 = ((~g26));
assign g11143 = (g10923&g4567);
assign II11477 = ((~g6488));
assign g10457 = ((~II15962));
assign II9581 = ((~g5111));
assign g2860 = ((~II5998));
assign g7470 = ((~g6927));
assign g11075 = ((~g10937));
assign II10367 = ((~g6234));
assign g7596 = ((~II12127))|((~II12128));
assign g5520 = ((~II8943));
assign II11122 = ((~g6450));
assign g6888 = ((~II10984));
assign g3708 = ((~II6867));
assign II12541 = ((~g7662));
assign II17528 = ((~g11487));
assign II11695 = ((~g7052));
assign II16496 = ((~g10707));
assign II13834 = ((~g8488));
assign g11480 = ((~g11456)&(~g4567));
assign g10380 = ((~II15864));
assign g7663 = ((~II12282));
assign g2531 = (g658&g668);
assign g3995 = ((~g3121));
assign g10591 = ((~II16258));
assign g2215 = ((~II5185))|((~II5186));
assign II14668 = ((~g9309));
assign g5248 = (g673&g4738);
assign g10700 = ((~II16379));
assign g2256 = ((~II5279));
assign g9534 = ((~II14687));
assign g7751 = ((~II12418));
assign g6695 = ((~II10666));
assign g7560 = ((~II12012));
assign g2219 = ((~g94));
assign II9287 = ((~g5576));
assign II14105 = ((~g8776));
assign g7772 = ((~II12481));
assign g4289 = ((~g4013));
assign II16066 = ((~g10428))|((~II16065));
assign g10251 = ((~g10195));
assign II5073 = ((~g34));
assign g6461 = ((~II10391));
assign g2022 = ((~g1346));
assign II16790 = ((~g10900));
assign g2987 = ((~g2481))|((~g883));
assign II12384 = ((~g7212));
assign II17546 = ((~g11500));
assign II14858 = (g9585)|(g9595)|(g9610)|(g9602);
assign g5033 = ((~II8406));
assign II12190 = ((~g7268));
assign g2338 = ((~g1909));
assign g3999 = (g1741&g2777);
assign g8421 = ((~II13577));
assign g4316 = (g1965&g3400);
assign II14242 = ((~g8787));
assign II11232 = ((~g6537));
assign g11041 = ((~II16784));
assign II14367 = ((~g8953));
assign II11704 = ((~g7008));
assign g3419 = ((~g3104));
assign II14257 = ((~g8805));
assign II9117 = ((~g5615));
assign II5343 = ((~g426))|((~II5341));
assign g7918 = ((~g7505));
assign II12300 = ((~g7240));
assign g2061 = ((~g1828));
assign II16024 = ((~g10426))|((~II16023));
assign II17277 = ((~g11390));
assign II16121 = ((~g10396));
assign g3097 = ((~g2482));
assign g8612 = ((~II13858))|((~II13859));
assign II5561 = ((~g869));
assign II10521 = ((~g822))|((~II10519));
assign g5500 = (g1657&g4272);
assign g11197 = ((~g11112));
assign g2538 = (g1466)|(g1458)|(II5649);
assign g7543 = ((~II11961));
assign II17255 = ((~g11344));
assign g7890 = ((~g7479));
assign g8290 = ((~II13224));
assign g5890 = ((~g5361));
assign g6707 = ((~g5949));
assign g2161 = (II5084&II5085);
assign g11176 = (g506&g11112);
assign II4883 = ((~g581));
assign II13876 = ((~g8535))|((~g1444));
assign g11291 = (g11247&g4233);
assign II13454 = ((~g8183));
assign g2556 = ((~g186));
assign g5708 = ((~II9253));
assign g6469 = (g5698)|(g4959);
assign II4987 = ((~g1003))|((~II4985));
assign g10642 = (g10612&g3829);
assign II14010 = ((~g8642));
assign g8214 = (g7472)|(g8004);
assign II15898 = ((~g857))|((~g10287));
assign g6639 = (g357&g6196);
assign g7465 = (g6876)|(g6410);
assign g3737 = ((~g2834));
assign g2331 = ((~g658));
assign g8655 = (g8532&g4013);
assign II12762 = ((~g7541));
assign g7823 = (g1923&g7479);
assign g6775 = (g822&g6231);
assign g5224 = (g4360)|(g3512);
assign II16586 = ((~g10850));
assign g6170 = ((~g5426));
assign g6116 = ((~II9801));
assign II8663 = ((~g4286))|((~II8662));
assign II7284 = ((~g3255));
assign g10101 = ((~II15335));
assign g8390 = (g8268&g6465);
assign g8377 = (g8185)|(g7958);
assign g11086 = ((~II16867));
assign g10890 = ((~II16632));
assign II12318 = ((~g6862));
assign II4973 = ((~g995))|((~II4971));
assign g8774 = (g5499)|(g8654);
assign g9747 = (g9173)|(g9509);
assign g5723 = ((~II9265));
assign II6714 = ((~g2961))|((~g201));
assign g5031 = (g1478&g4640);
assign g11347 = ((~II17164));
assign g7792 = ((~II12541));
assign g8737 = ((~g2317))|((~g4921))|((~g8688));
assign g10850 = ((~II16550));
assign g4263 = ((~g3586));
assign g4336 = ((~g4130));
assign g5509 = ((~g4739));
assign g8966 = (g8081&g6778&g8849);
assign II10759 = ((~g5803));
assign II15296 = ((~g9995));
assign g6324 = (g1240&g5949);
assign g4426 = ((~g3914));
assign g3625 = ((~II6771))|((~II6772));
assign g2131 = ((~II5060));
assign g4912 = ((~II8282));
assign II11085 = ((~g6433));
assign g9415 = (g1733&g9052);
assign II14239 = ((~g8803));
assign g9720 = (g1546&g9490);
assign II5626 = (g521)|(g525)|(g530)|(g534);
assign II17213 = ((~g11290));
assign II5284 = ((~g762))|((~II5282));
assign g7540 = ((~II11956));
assign g9845 = ((~g9679));
assign g7259 = ((~II11494));
assign g4081 = ((~II7210));
assign II11942 = ((~g6909));
assign g3907 = ((~II7076));
assign g10425 = ((~g10293)&(~g4620));
assign II7946 = ((~g3417));
assign g6127 = ((~II9826));
assign II16604 = ((~g10786));
assign II7396 = ((~g4102));
assign g10549 = (g4951)|(g10451);
assign II6074 = ((~g2228));
assign g4538 = ((~g3475))|((~g2399));
assign g4788 = (g511&g3436);
assign g5094 = ((~II8462));
assign g5263 = (g709&g4761);
assign II10952 = ((~g6556));
assign g7184 = (g6625)|(g6047);
assign II6504 = ((~g3214));
assign II6233 = ((~g2299));
assign g3460 = ((~II6665))|((~II6666));
assign g5241 = ((~g4386));
assign g4514 = ((~g3946));
assign II10932 = ((~g5555))|((~II10930));
assign g11278 = (g11253)|(g11150);
assign II12589 = ((~g7571));
assign g5825 = (g3204&g5318);
assign g9192 = (g6454&g8955);
assign II11420 = ((~g6417));
assign II8506 = ((~g4334));
assign II11653 = ((~g6954));
assign II8123 = ((~g3630));
assign g10190 = ((~II15548));
assign II17302 = ((~g11391));
assign II11936 = ((~g7004))|((~II11935));
assign II6947 = ((~g2860));
assign g11148 = (g2321&g10913);
assign g3813 = ((~II7034))|((~II7035));
assign g4592 = ((~g3829));
assign g3812 = ((~g3228));
assign g7303 = (g7145)|(g6329);
assign g11539 = ((~g11519));
assign II15338 = ((~g10013));
assign g9025 = ((~II14412));
assign g11320 = (g11201&g4379);
assign g11416 = ((~II17296))|((~II17297));
assign II14204 = ((~g591))|((~II14202));
assign g10056 = ((~II15275));
assign g4250 = ((~g3698));
assign II11049 = ((~g6635));
assign g8626 = ((~g8498));
assign g2644 = ((~g1990));
assign g6802 = ((~II10816));
assign II16214 = ((~g10500));
assign g4521 = ((~g3586));
assign g9698 = (g1571&g9474);
assign g8173 = (g7971&g3112);
assign II12499 = ((~g7725));
assign II10706 = ((~g6080));
assign II7729 = ((~g3757));
assign g9782 = ((~II14933));
assign g8336 = ((~II13388));
assign g8331 = ((~II13373));
assign g6038 = (g5528)|(g3979);
assign II8640 = ((~g4278))|((~g516));
assign g6288 = ((~II10123));
assign II6789 = ((~g2748));
assign g1965 = ((~g119));
assign g3545 = ((~II6733));
assign g9519 = (g9173)|(g9151)|(g9125);
assign II12056 = ((~g6929));
assign II7659 = ((~g3731));
assign II13445 = ((~g8149));
assign g11637 = (g11626&g5446);
assign g10799 = (g6225)|(g10769);
assign II15694 = ((~g10234));
assign II14678 = ((~g9265));
assign II5070 = ((~g1194));
assign II7118 = ((~g2979));
assign II13258 = ((~g1900))|((~g8153));
assign g10051 = ((~II15272));
assign g4217 = ((~II7468));
assign g3753 = ((~g2382))|((~g2364))|((~g2800));
assign g6624 = (g348&g6171);
assign g11265 = (g11189)|(g11027);
assign g9703 = (g1577&g9474);
assign g6315 = ((~II10204));
assign g5886 = ((~g5361));
assign II13952 = ((~g8451));
assign II10861 = ((~g6694));
assign II8324 = ((~g4794));
assign g5639 = ((~II9080));
assign g3940 = ((~g2920));
assign g8236 = (g7526)|(g8001);
assign II12223 = ((~g7049));
assign g5482 = ((~II8903));
assign II9776 = ((~g5353));
assign g7438 = ((~g7232));
assign II16676 = ((~g10798));
assign g5569 = (g4816&g2338);
assign g5107 = ((~g4459));
assign g7334 = ((~II11650));
assign g3942 = (g219&g3164);
assign II13489 = ((~g8233));
assign g3967 = ((~g3247));
assign II14119 = ((~g8779));
assign II5516 = ((~g1260))|((~g1019));
assign g6019 = ((~g617))|((~g4921));
assign g8359 = ((~II13457));
assign g10169 = ((~II15503));
assign g2825 = ((~II5935));
assign II9857 = ((~g5269));
assign g11605 = (g11584)|(g11555);
assign g8416 = (g731&g8151);
assign g3520 = ((~g2779));
assign g11209 = (g11074&g9448);
assign g4766 = ((~g3440));
assign g6443 = ((~g6157));
assign II4966 = ((~g330))|((~II4964));
assign g9725 = (g9642)|(g9659)|(g9616)|(II14862);
assign g11646 = ((~II17742));
assign II14217 = ((~g8826))|((~II14216));
assign II5410 = ((~g901));
assign g3978 = ((~g3207))|((~g1822));
assign g8451 = (g3440)|(g8366);
assign g6582 = ((~g5949));
assign g6432 = ((~g6146));
assign g4739 = ((~g4117));
assign g11309 = ((~II17096));
assign II9433 = ((~g5069));
assign g4878 = (g1868&g3531);
assign g6904 = ((~II11008));
assign g9813 = ((~II14948));
assign g5917 = (g1044&g5320);
assign g10244 = ((~g10131));
assign g4113 = ((~II7255));
assign g11229 = (g11154)|(g11012);
assign g8147 = (g2955&g7961);
assign II5311 = ((~g98));
assign II12159 = ((~g7243));
assign g10579 = ((~g10528));
assign g4339 = ((~g4144));
assign g6964 = ((~g6509));
assign II13354 = ((~g8214));
assign g6560 = ((~g5759));
assign II17265 = ((~g11352));
assign g8439 = ((~II13615));
assign g5116 = ((~g4682));
assign g9642 = (g2654&g9240);
assign g2623 = ((~g1999));
assign II12793 = ((~g7619));
assign II8911 = ((~g4565));
assign g10886 = ((~g10807))|((~g10805));
assign II14531 = ((~g9273));
assign g10658 = (g10595)|(g7674);
assign II15870 = ((~g10358))|((~g2713));
assign g10932 = ((~g10827));
assign g8195 = ((~II13122));
assign II13990 = ((~g622))|((~g8688));
assign g10121 = ((~II15371));
assign II14970 = ((~g9732));
assign g2176 = ((~g82));
assign II7636 = ((~g3330));
assign g9658 = (g947&g9240);
assign g4141 = (g2707&g3051);
assign II11632 = ((~g6931));
assign II6805 = ((~g3268))|((~g471));
assign g2507 = ((~II5584));
assign g11475 = ((~II17466));
assign g2890 = ((~II6052));
assign g9966 = (g9956&g9536);
assign II8024 = ((~g4117));
assign g9864 = (g1604&g9778);
assign II6510 = ((~g3267));
assign II4954 = ((~g401))|((~g327));
assign II14485 = ((~g8883));
assign g8089 = ((~g7934));
assign II12627 = ((~g7697));
assign g7929 = ((~g7519));
assign g4050 = ((~II7163));
assign g10317 = ((~II15749));
assign g5416 = ((~II8851));
assign II9575 = ((~g5608))|((~II9574));
assign II5605 = ((~g1149))|((~II5604));
assign g3790 = ((~g3228));
assign g6875 = (g1905&g6400);
assign II13285 = ((~g8159))|((~II13283));
assign g8514 = ((~II13711));
assign g9803 = ((~g9392)&(~g9367));
assign g8265 = (g7881)|(g3396);
assign g7574 = ((~g6995));
assign II16799 = ((~g11017));
assign g11463 = (g11432&g5446);
assign g2854 = ((~II5986));
assign g11288 = (g11204)|(g11070);
assign g11212 = (g944&g11155);
assign g11152 = (g369&g10903);
assign II17318 = ((~g11340));
assign g6341 = (g272&g5885);
assign g11096 = ((~II16879));
assign g10432 = ((~g10350)&(~g3566));
assign II15193 = ((~g9968));
assign g5299 = ((~g4393));
assign II13017 = ((~g7848));
assign g10676 = ((~g10570));
assign II17552 = ((~g11502));
assign g10876 = ((~II16598));
assign II10927 = ((~g6755));
assign II16638 = ((~g10863));
assign g4893 = (g635&g4739);
assign II12282 = ((~g7113));
assign g5677 = ((~II9188));
assign II12838 = ((~g7682));
assign II8253 = ((~g4637));
assign g8284 = (g8102)|(g7821);
assign g6274 = ((~II10081));
assign g7232 = ((~II11472));
assign g6247 = (g127&g5361);
assign II11566 = ((~g6820));
assign g6728 = (g6250&g4318);
assign II5893 = ((~g2057))|((~II5891));
assign g9817 = ((~g9392)&(~g9367));
assign g5100 = (g1791&g4606);
assign g1975 = ((~g622));
assign II6220 = ((~g883));
assign g5182 = (g1240&g4713);
assign g7692 = ((~g7148));
assign II15209 = (g8169)|(g9905)|(g9934)|(g9830);
assign g5731 = (g1583&g5175);
assign II10607 = ((~g5763));
assign g6816 = ((~II10858));
assign g8127 = (g1927&g7949);
assign g10087 = ((~II15314));
assign II11686 = ((~g7039));
assign g11097 = (g378&g10884);
assign II11094 = ((~g6657));
assign g8812 = (g7939)|(g8724);
assign g7651 = (g7135)|(g4084);
assign II13245 = ((~g8269));
assign II6356 = ((~g2459));
assign II8848 = ((~g4490));
assign g4934 = ((~g4243));
assign II9141 = ((~g5402));
assign II6580 = ((~g3186));
assign g5613 = ((~g4840));
assign g2344 = ((~II5410));
assign II7820 = ((~g3811));
assign II4929 = ((~g391))|((~II4928));
assign g8649 = (g8499)|(g4519);
assign II8717 = ((~g4052))|((~II8715));
assign II11800 = ((~g7246));
assign g2270 = ((~II5311));
assign II11975 = ((~g1462))|((~II11973));
assign g8729 = ((~g8595));
assign g4490 = (g1141&g3913);
assign g5841 = (g4914)|(g4230);
assign g2677 = ((~g2034));
assign II8228 = ((~g4468));
assign g3037 = ((~g2135));
assign g5029 = (g1077&g4521);
assign g10974 = ((~II16723));
assign g9838 = (g9700&g9754);
assign g4499 = ((~g3546));
assign g2940 = (g2424&g1654);
assign g3246 = ((~g2482));
assign II16196 = ((~g10496));
assign II10201 = ((~g5998));
assign g8979 = ((~II14358));
assign g7619 = ((~II12205));
assign g3860 = (g3107)|(g2167);
assign II6080 = ((~g2108));
assign II11348 = ((~g6695));
assign g3112 = ((~g2482));
assign g10735 = ((~II16416));
assign II13320 = ((~g8096));
assign g9613 = (g1176&g9125);
assign g6832 = (g1383&g6596);
assign g11654 = ((~II17764));
assign g4272 = ((~g3586));
assign II5438 = ((~g18));
assign II12400 = ((~g7537));
assign II12032 = ((~g6923));
assign g6031 = ((~II9642));
assign g5772 = (g1555&g5214);
assign g10138 = ((~II15412));
assign II11537 = ((~g7144));
assign II14709 = ((~g9267));
assign g7519 = ((~g6956));
assign g10439 = ((~g10334));
assign II13645 = ((~g8379));
assign II16200 = ((~g10494));
assign g5189 = (g4345)|(g3496);
assign II15190 = ((~g9974));
assign g8730 = (g8613&g7917);
assign II17733 = ((~g11639));
assign g3938 = ((~g2991));
assign g5818 = ((~g5320));
assign II15526 = ((~g10051));
assign II12062 = ((~g1478))|((~II12060));
assign g4671 = ((~g3354));
assign g5286 = ((~II8751))|((~II8752));
assign g2056 = ((~II4859));
assign g7780 = ((~II12505));
assign II17500 = ((~g11478));
assign g4820 = (g186&g3946);
assign II11790 = ((~g7246));
assign II14444 = ((~g1834))|((~II14442));
assign II6976 = ((~g2884));
assign g8878 = (g8099&g6368&g8858);
assign II12412 = ((~g7520));
assign II6676 = ((~g2759));
assign II9525 = ((~g5001));
assign g10401 = (g9317)|(g10291);
assign g2500 = ((~g178))|((~g182));
assign g11433 = ((~II17350));
assign g4827 = (g213&g3946);
assign g8868 = ((~II14176));
assign g11220 = (g962&g11054);
assign g10540 = ((~II16187));
assign II13918 = ((~g8451));
assign g8109 = ((~g5052))|((~g7853));
assign II12430 = ((~g7649));
assign g6296 = ((~II10147));
assign g7846 = (g7722)|(g7241);
assign II12409 = ((~g7501));
assign g7009 = ((~II11152));
assign II4948 = ((~g586));
assign II9620 = ((~g5189));
assign g11028 = (g396&g10974);
assign II5658 = ((~g560));
assign g3878 = ((~g2920));
assign g2757 = ((~II5837));
assign II13618 = ((~g8345));
assign II9171 = ((~g4902));
assign g5719 = ((~II9259));
assign g6846 = ((~II10910));
assign II9965 = ((~g5493));
assign g8329 = ((~II13367));
assign g3758 = ((~II6955));
assign g8505 = (g8309&g4789);
assign II6111 = ((~g1494))|((~II6109));
assign g2945 = (g2411&g1684);
assign g2611 = ((~II5734));
assign g6137 = ((~II9848));
assign g8708 = (g7605&g8592);
assign g2046 = ((~g1845));
assign g9828 = (g9722&g9785);
assign II17158 = ((~g11312));
assign g6347 = (g275&g5890);
assign II13370 = ((~g8128));
assign II16458 = ((~g10734));
assign g10080 = ((~II15308));
assign g6003 = ((~g5552))|((~g5548));
assign II11590 = ((~g6829));
assign g10564 = (g10560)|(g7368);
assign II11677 = ((~g7056));
assign g10234 = ((~g10188));
assign g6412 = ((~II10322));
assign g6485 = (g5848)|(g5067);
assign g6385 = ((~g6119));
assign g9593 = (g898&g9205);
assign g3705 = ((~g3113));
assign II9105 = ((~g5589));
assign II8625 = ((~g4267))|((~II8624));
assign g11496 = ((~II17504))|((~II17505));
assign g8934 = ((~II14278))|((~II14279));
assign II13504 = ((~g677))|((~g8247));
assign g5314 = ((~g4387));
assign g6332 = (g1374&g5904);
assign II5388 = ((~g889));
assign II8237 = ((~g4295));
assign II15617 = ((~g10153))|((~II15615));
assign g4887 = ((~II8234));
assign g9911 = (g9846)|(g9689);
assign g3207 = ((~g2439));
assign II8462 = ((~g4475));
assign g8003 = ((~II12835));
assign g7573 = ((~II12046))|((~II12047));
assign g8140 = ((~II13017));
assign g10478 = ((~II16052))|((~II16053));
assign g8157 = (g7965)|(g7623);
assign II5366 = (g1280)|(g1284)|(g1292)|(g1296);
assign II15320 = ((~g10013));
assign g7581 = (g7092&g5420);
assign g7532 = ((~II11932));
assign g4713 = ((~g3546));
assign II6661 = ((~g2752));
assign g7443 = ((~II11841));
assign g9413 = ((~II14613))|((~II14614));
assign g2911 = (g2411&g1675);
assign g5145 = (g1639&g4673);
assign g9661 = ((~II14786));
assign II6520 = ((~g3186));
assign g5811 = ((~II9415));
assign II10018 = ((~g5862));
assign g11413 = (g11354&g10679);
assign g7510 = (g7186)|(g6730);
assign II7763 = ((~g3769));
assign g7189 = (g6632)|(g6053);
assign g10865 = (g5538)|(g10752);
assign g8560 = ((~II13773));
assign g11150 = (g3087&g10913);
assign g6145 = ((~II9860));
assign g7584 = ((~II12075))|((~II12076));
assign g10745 = (g10658&g3586);
assign g7966 = ((~II12762));
assign g4465 = (g1117&g3828);
assign g7394 = ((~II11778));
assign g5664 = ((~II9153));
assign g6122 = (g5172)|(g5180);
assign g8014 = (g7740&g7419);
assign g7959 = ((~II12751));
assign g3723 = ((~g3071));
assign II7300 = ((~g2883));
assign g4164 = ((~II7311));
assign II12577 = ((~g7532));
assign g8254 = (g2773&g7909);
assign II9557 = ((~g5598))|((~g782));
assign g8881 = ((~II14210))|((~II14211));
assign II9947 = ((~g5233))|((~II9946));
assign g10696 = ((~g10621));
assign g9995 = (II15199)|(II15200);
assign II13806 = ((~g8478));
assign g5779 = ((~II9371));
assign g11107 = ((~g10974));
assign g8274 = ((~II13194));
assign g8267 = (g7889)|(g3422);
assign g3799 = ((~II7022));
assign g5934 = (g5215&g1965);
assign II7438 = ((~g3461));
assign II11011 = ((~g6340));
assign g9734 = (g9415)|(g9428)|(g9421);
assign g10325 = (g10248&g3307);
assign g6546 = (g5796)|(g5026);
assign g10670 = (g10571&g9091);
assign g8297 = ((~II13245));
assign g7631 = ((~II12235));
assign g6733 = (g5678&g4324);
assign g3389 = (g207&g3228);
assign g6758 = ((~II10770))|((~II10771));
assign g3011 = ((~g591))|((~g2382));
assign g6531 = (g79&g6056);
assign g7767 = ((~II12466));
assign g2316 = (g1300)|(g1304)|(g1270)|(II5366);
assign g9586 = (g2727&g9173);
assign g3719 = ((~g2920));
assign II5468 = ((~g1245))|((~g999));
assign II10739 = ((~g5942));
assign g8388 = (g8177&g7689);
assign II16817 = ((~g10912));
assign g2006 = ((~g932));
assign II8575 = ((~g4234))|((~g496));
assign g8839 = ((~g8750))|((~g4401));
assign g7853 = ((~II12652));
assign g8697 = ((~g8660));
assign g8150 = ((~II13039));
assign g7886 = ((~g7479));
assign g7256 = ((~II11489));
assign g4174 = ((~II7339));
assign II4912 = ((~g318))|((~II4910));
assign g8552 = (g8217)|(g8388);
assign II9851 = ((~g5405));
assign g7502 = ((~II11882));
assign g10452 = (g10439&g3388);
assign II16073 = ((~g845))|((~II16072));
assign g8714 = ((~II14005));
assign II10630 = ((~g5889));
assign g6306 = ((~II10177));
assign g7293 = (g7063)|(g6319);
assign g10433 = ((~g10330)&(~g3507));
assign g2872 = ((~II6016));
assign II9839 = ((~g5226));
assign g11435 = ((~II17356));
assign g6709 = ((~g5949));
assign II7509 = ((~g3566));
assign II9213 = ((~g4944));
assign g2506 = ((~g636));
assign g2350 = ((~II5424));
assign g6580 = (g1801&g5944);
assign II8315 = ((~g4788));
assign g10818 = (g10730&g4545);
assign g4013 = ((~II7157));
assign g2227 = ((~g95));
assign g2209 = ((~g93));
assign II14443 = ((~g8970))|((~II14442));
assign g10063 = ((~II15287));
assign g11404 = ((~II17255));
assign g7741 = (g6961&g3880);
assign II9845 = ((~g5405));
assign II6914 = ((~g2828));
assign g7722 = (g7127&g6449);
assign II11450 = ((~g6488));
assign g10392 = ((~II15891))|((~II15892));
assign II10843 = ((~g6723));
assign g5174 = (g1235&g4681);
assign g11452 = ((~II17413));
assign g11443 = (g7130)|(g11407);
assign g4905 = (g1853&g4243);
assign II11935 = ((~g7004))|((~g1458));
assign g4906 = ((~II8275));
assign II12136 = ((~g7110))|((~g131));
assign g6826 = (g225&g6596);
assign g5859 = ((~g3362)&(~g4943));
assign II9377 = ((~g5576));
assign g8573 = ((~II13812));
assign g6318 = (g1300&g5949);
assign g4993 = (g1448&g4682);
assign g7697 = ((~g7101));
assign g4463 = ((~g3829));
assign g10075 = ((~II15302));
assign II11970 = ((~g6918));
assign g6337 = ((~II10234));
assign II7668 = ((~g3733));
assign II5221 = ((~g1407));
assign g3776 = ((~g2579));
assign g9856 = (g1592&g9773);
assign g10860 = (g5513)|(g10743);
assign II15048 = (g7853)|(g9683)|(g9624)|(g9785);
assign g10628 = ((~II16307));
assign g11203 = ((~g11112));
assign g4298 = ((~g4130));
assign II14561 = ((~g9025));
assign g8635 = ((~II13918));
assign g4541 = ((~II7946));
assign g8828 = ((~g8744));
assign II10620 = ((~g5884));
assign II9224 = ((~g5063));
assign II17410 = ((~g11419));
assign g3041 = ((~g2364))|((~g2399))|((~g2374))|((~g2382));
assign g8234 = ((~g7826));
assign g6912 = (g6350)|(g4235);
assign II6287 = ((~g2091))|((~g981));
assign g7374 = ((~II11752));
assign g5121 = ((~g4682));
assign g6515 = (g5739)|(g4993);
assign II6447 = ((~g2264))|((~g1776));
assign g9427 = ((~g9079));
assign g7710 = (g700&g7214);
assign g7050 = (g5896&g6575);
assign g11579 = (g5123)|(g11551);
assign g2763 = ((~II5847));
assign g10032 = ((~II15232));
assign g5839 = ((~II9452));
assign II14546 = ((~g9312));
assign g11183 = ((~II16950));
assign g7076 = ((~II11303));
assign II14249 = ((~g8804));
assign g10682 = (g10600&g3863);
assign g3373 = ((~II6565));
assign g6425 = ((~g6141));
assign g4003 = ((~g3144));
assign g8180 = ((~II13090))|((~II13091));
assign g8379 = ((~II13485));
assign g5643 = ((~II9090));
assign g11244 = ((~g11112));
assign II9519 = ((~g4998));
assign II7766 = ((~g3770));
assign g6854 = ((~II10920));
assign g4762 = ((~II8116));
assign g8694 = ((~II13975));
assign g8272 = ((~II13188));
assign g10305 = ((~II15725));
assign g10227 = ((~II15601));
assign II16298 = ((~g10553));
assign g11380 = (g11321&g4285);
assign g11627 = ((~II17695));
assign II5579 = ((~g1197));
assign g11582 = (g1311&g11540);
assign II17170 = ((~g11294));
assign II9923 = ((~g5308));
assign II9602 = ((~g5013));
assign g6724 = ((~II10719));
assign g7287 = ((~II11537));
assign g8252 = (g7988)|(g7679);
assign g5592 = ((~II9007))|((~II9008));
assign g7909 = ((~g7664));
assign g3717 = ((~II6880))|((~II6881));
assign g10867 = ((~II16571));
assign g3988 = ((~g3121));
assign II11021 = ((~g6398));
assign g4785 = ((~g3337));
assign II6747 = ((~g2938))|((~II6746));
assign II6837 = ((~g3287))|((~II6836));
assign II8234 = ((~g4232));
assign II6778 = ((~g2892))|((~II6777));
assign g6927 = ((~II11049));
assign II17179 = ((~g11307));
assign g2322 = ((~II5378));
assign g10359 = ((~g10227)&(~g4620));
assign g5751 = ((~II9323));
assign g7125 = (g1212&g6648);
assign g6787 = (g266&g5875);
assign g3392 = ((~g3121));
assign g5903 = ((~II9536));
assign g10718 = (g6238)|(g10706);
assign g7033 = ((~II11188));
assign II7333 = ((~g3729));
assign II6624 = ((~g2629));
assign II9860 = ((~g5405));
assign g10574 = ((~II16239));
assign g4172 = ((~II7333));
assign g7368 = (g6980&g3880);
assign II11249 = ((~g6541));
assign II6091 = ((~g2270));
assign II11278 = ((~g305))|((~g6485));
assign g4746 = ((~II8098));
assign II10012 = ((~g5543));
assign II8080 = ((~g3538));
assign g9555 = (g9107&g3391);
assign g2903 = ((~g2166));
assign g9088 = (g8927)|(g8381);
assign gbuf11 = (g1206);
assign II10756 = ((~g5810));
assign g4486 = (g1711&g3910);
assign g2814 = ((~II5916));
assign g5735 = ((~II9293));
assign g10635 = (g10622)|(g7732);
assign II5837 = ((~g2507));
assign g6407 = ((~II10317));
assign II6144 = ((~g1976))|((~II6143));
assign g8060 = (g7593&g5919);
assign g7361 = ((~II11731));
assign II17356 = ((~g11384));
assign g8043 = (g7582&g5128);
assign g11415 = ((~II17289))|((~II17290));
assign g6166 = ((~II9893));
assign g7265 = (g6756)|(g6204);
assign II5805 = (g2102)|(g2099)|(g2096)|(g2088);
assign g5510 = (g1630&g4280);
assign II9394 = ((~g5195));
assign g3424 = ((~g2896));
assign g2034 = ((~g1766));
assign II8011 = ((~g3820));
assign g4203 = ((~II7426));
assign II8490 = ((~g4526));
assign g2517 = ((~II5619))|((~II5620));
assign g5118 = ((~g2439))|((~g4806))|((~g4073));
assign II17435 = ((~g11454));
assign g6906 = (g6791)|(g5674);
assign II12638 = ((~g7708));
assign g4270 = ((~g4013));
assign II14077 = ((~g8758));
assign g4185 = ((~II7372));
assign g2877 = ((~II6025));
assign g2510 = ((~II5592))|((~II5593));
assign g8873 = ((~II14191));
assign g8184 = ((~II13105));
assign II17441 = ((~g11445));
assign g2238 = ((~II5237));
assign g11372 = (g11316&g4266);
assign g6834 = (g1365&g6596);
assign II11540 = ((~g6877));
assign g2799 = ((~g2276));
assign g7961 = ((~g7664));
assign g10290 = ((~II15694));
assign II11810 = ((~g7246));
assign II10503 = ((~g5858));
assign g11279 = (g4939&g11200);
assign II10682 = ((~g6051));
assign g7353 = ((~II11707));
assign g1994 = ((~g794));
assign II7351 = ((~g4061));
assign II8139 = ((~g3681));
assign g2804 = (g2132&g1891);
assign g8794 = ((~II14109));
assign g5205 = ((~g4366));
assign g4582 = (g525&g4055);
assign II5677 = ((~g1223))|((~II5675));
assign II14499 = ((~g8889));
assign g9617 = (g9&g9274);
assign g6105 = (g5279)|(g4559);
assign g4577 = ((~II7984));
assign g11281 = (g4948&g11202);
assign g5398 = (g4610&g2224);
assign II13039 = ((~g8054));
assign II6880 = ((~g3301))|((~II6879));
assign g6058 = (g1035&g5320);
assign g9897 = (g9884&g9624);
assign II12610 = ((~g7627));
assign g8786 = (g8638&g8716);
assign g2234 = ((~g87));
assign II5127 = ((~g1386))|((~II5126));
assign g4476 = ((~g3807))|((~g3071));
assign g9957 = (g9949)|(g9943)|(g9776);
assign II15308 = ((~g10019));
assign g7920 = ((~g7516));
assign g11598 = ((~II17642));
assign g11459 = (g11427&g5446);
assign g11393 = (g11280&g7916);
assign g2121 = ((~II5041));
assign II13439 = ((~g8187));
assign g9312 = ((~II14509));
assign g7346 = ((~II11686));
assign g10261 = ((~g10126));
assign g2269 = ((~II5308));
assign g6448 = ((~II10374));
assign II15269 = ((~g9993));
assign II8499 = ((~g4330));
assign g2896 = ((~g2356));
assign g10424 = ((~g10292)&(~g4620));
assign II9323 = ((~g5620));
assign II10258 = ((~g6134));
assign g10207 = ((~g10186));
assign g7459 = (g7148&g2814);
assign g11055 = ((~g10950));
assign II11898 = ((~g6896));
assign g5523 = (g1663&g4290);
assign II5649 = (g1499)|(g1486)|(g1482);
assign g5620 = ((~g4417));
assign g8322 = (g8136)|(g6891);
assign g8345 = ((~II13415));
assign II16667 = ((~g10780));
assign g3271 = ((~II6443));
assign g8745 = ((~g8617))|((~g6517))|((~g6964));
assign g10554 = (g4097)|(g10503);
assign g5851 = (g4941)|(g4253);
assign g5742 = ((~II9308));
assign g10899 = ((~g10803));
assign g5502 = (g1932&g4275);
assign g7036 = ((~g6420));
assign II5263 = ((~g456))|((~g461));
assign II8278 = ((~g4495));
assign g5027 = ((~II8396));
assign II17739 = ((~g11641));
assign g2557 = ((~g1840));
assign g4590 = ((~II7999));
assign II5599 = (g516)|(g511)|(g506)|(g501);
assign g5705 = ((~II9248));
assign g5808 = ((~g5320));
assign II16169 = ((~g10448));
assign g5091 = ((~g4385));
assign g8810 = (g7933)|(g8720);
assign g7927 = ((~g7500));
assign g5651 = ((~II9114));
assign II11100 = ((~g6442));
assign g6573 = ((~II10508))|((~II10509));
assign g3664 = ((~g3209));
assign g3500 = ((~II6690));
assign g9891 = (g9741)|(g9760);
assign II17206 = ((~g11323));
assign II7456 = ((~g3716));
assign II9956 = ((~g5485));
assign g11065 = ((~g10974));
assign II16484 = ((~g10770));
assign II9505 = ((~g5088));
assign g5800 = ((~II9402));
assign g8476 = ((~II13674));
assign g9922 = (g9864)|(g9705);
assign II11269 = ((~g6545));
assign II12286 = ((~g7231));
assign g2792 = ((~II5879))|((~II5880));
assign g4533 = ((~II7938));
assign g9929 = (g9871)|(g9718);
assign g9390 = (g1333&g9151);
assign g7719 = (g718&g7227);
assign g6919 = ((~g6453));
assign II5041 = ((~g1179));
assign g6430 = (g5044&g5791);
assign g11397 = ((~II17234));
assign II6143 = ((~g1976))|((~g646));
assign II16500 = ((~g10711));
assign II13128 = ((~g7976));
assign g4255 = (g4009)|(g4047);
assign II5963 = ((~g2179));
assign II6317 = (g2406&g2420&g2434&g2438);
assign II5427 = ((~g913));
assign g6557 = ((~g5748));
assign II15583 = ((~g10157));
assign g9591 = ((~g9125)&(~g9151));
assign g11591 = (g2988&g11561);
assign II16610 = ((~g10792));
assign g7599 = ((~II12144))|((~II12145));
assign g8305 = ((~II13284))|((~II13285));
assign g7607 = ((~II12171));
assign g2750 = ((~II5818));
assign g5683 = ((~II9202));
assign g4950 = (g1415&g4682);
assign g6584 = ((~II10538));
assign g4348 = (g3497&g1909);
assign g3543 = ((~g3101));
assign g6503 = ((~II10421));
assign II12683 = ((~g7387));
assign g11329 = (g11302)|(g11169);
assign g6041 = ((~II9658));
assign II13206 = ((~g8197));
assign II5164 = ((~g1508))|((~g1499));
assign g11589 = (g1333&g11548);
assign g10855 = (g6075)|(g10736);
assign II11725 = ((~g7040));
assign II8851 = ((~g4498));
assign g8406 = (g695&g8131);
assign g6793 = ((~II10795));
assign g6949 = ((~II11091));
assign g4415 = ((~g3914));
assign g11012 = (g5196&g10827);
assign II10984 = ((~g6757));
assign g4988 = ((~II8358));
assign g10441 = ((~g10351)&(~g3566));
assign II15749 = ((~g10263));
assign II7642 = ((~g3440));
assign g4605 = ((~g3077)&(~g2669)&(~g3485)&(~g2655));
assign g10289 = ((~II15691));
assign II17657 = ((~g11598));
assign g3431 = (g2951)|(g2957);
assign g4831 = (g810&g4109);
assign g4070 = (g3263&g2330);
assign II15891 = ((~g853))|((~II15890));
assign g2005 = ((~g928));
assign g10822 = ((~II16534));
assign II8476 = ((~g4577));
assign II7151 = ((~g2642));
assign g8535 = ((~II13744));
assign II10096 = ((~g5794));
assign II12783 = ((~g7590));
assign II9935 = ((~g5477));
assign II16280 = ((~g10537));
assign II10846 = ((~g6729));
assign g6282 = ((~II10105));
assign g3531 = ((~g2971));
assign II10828 = ((~g6708));
assign g2957 = (g2424&g1663);
assign g10367 = (g10362&g3375);
assign g4589 = ((~II7996));
assign g9823 = ((~II14970));
assign g9762 = ((~II14903));
assign g6641 = ((~II10598));
assign g7898 = (g7511&g7041);
assign II9486 = ((~g5066));
assign g10162 = ((~II15482));
assign g6920 = ((~II11034));
assign g10884 = ((~g10809));
assign g9886 = (g9607)|(g9592)|(g9759);
assign g6051 = ((~II9680));
assign g8827 = (g8552&g8696);
assign g10556 = (g4115)|(g10506);
assign II7176 = ((~g2623));
assign g5213 = ((~g4640));
assign II6193 = ((~g2155));
assign g2336 = ((~g1900));
assign g8958 = ((~II14323));
assign g6932 = ((~II11058));
assign g11603 = (g11582)|(g11553);
assign g2107 = ((~II4986))|((~II4987));
assign g7349 = ((~II11695));
assign g4184 = ((~II7369));
assign g5567 = ((~II8982));
assign g10170 = ((~g10118));
assign g9905 = (g9872&g9680);
assign g8843 = ((~g8542))|((~g8757))|((~g8545));
assign g6565 = ((~g5790));
assign g11353 = ((~II17176));
assign g8980 = ((~II14361));
assign II17713 = ((~g11621));
assign g4383 = (g2517&g3829);
assign g5879 = ((~II9498));
assign g8723 = ((~g8585));
assign II5619 = ((~g1766))|((~II5618));
assign II17070 = ((~g11233));
assign g4718 = (g650&g3343);
assign g10280 = ((~g10160));
assign g4293 = (g4064)|(g4068);
assign g5267 = ((~II8711));
assign II11608 = ((~g6903));
assign II17234 = ((~g11353));
assign g11019 = (g421&g10974);
assign g10910 = ((~II16682));
assign II7157 = ((~g3015));
assign g7776 = ((~II12493));
assign g8414 = ((~II13553))|((~II13554));
assign g11225 = (g11149)|(g11009);
assign g6264 = ((~II10051));
assign II6726 = ((~g3306));
assign II13317 = ((~g8093));
assign II9090 = ((~g5567));
assign II16660 = ((~g10793));
assign II14558 = ((~g9024));
assign g3363 = ((~II6549));
assign g5686 = (g158&g5361);
assign g7948 = (g2855&g7497);
assign II17584 = ((~g11354))|((~g11515));
assign g7206 = ((~II11436));
assign g2100 = ((~II4948));
assign g2979 = ((~II6208))|((~II6209));
assign g8763 = (g7440&g8680);
assign II15326 = ((~g10025));
assign g4522 = (g360&g3586);
assign g7337 = ((~II11659));
assign g11428 = ((~II17337));
assign g6861 = ((~II10941));
assign II12045 = ((~g6951))|((~g1486));
assign g6204 = (g3738&g4921);
assign g10372 = ((~g10345)&(~g3463));
assign II9883 = ((~g5557));
assign g2431 = ((~II5510));
assign II6955 = ((~g2871));
assign g6971 = ((~g6517));
assign II10111 = ((~g5754));
assign g6894 = (g6763)|(g4868);
assign g8318 = ((~II13338));
assign g5669 = ((~II9168));
assign g6868 = ((~II10946));
assign g3164 = ((~II6370));
assign g5221 = (g1260&g4730);
assign g5273 = (g1074&g4776);
assign g6939 = ((~II11071));
assign g4614 = ((~g3829));
assign II17678 = ((~g11607));
assign g10768 = (g10649&g4840);
assign II7372 = ((~g4057));
assign g11625 = (g6535)|(g11597);
assign g8606 = ((~g8481));
assign II10434 = ((~g5843));
assign II10698 = ((~g5856));
assign g5999 = ((~g2753)&(~g4953));
assign g8441 = ((~II13621));
assign g10906 = ((~II16670));
assign g9654 = ((~g9125)&(~g9173));
assign g9691 = (g269&g9432);
assign II13539 = ((~g8157))|((~II13537));
assign g6177 = (g5444)|(g4712);
assign II10795 = ((~g6123));
assign g10345 = ((~II15801));
assign g4370 = ((~II7671));
assign g9557 = (g9052)|(g9030);
assign g1997 = ((~g798));
assign g10362 = ((~g10228)&(~g3507));
assign g6688 = ((~II10655));
assign g10620 = ((~II16295));
assign g6131 = ((~g5548));
assign g7931 = (g2809&g7446);
assign g4555 = ((~II7964));
assign II12559 = ((~g7477));
assign g10787 = ((~II16487));
assign g7527 = ((~g7148));
assign g6097 = ((~II9754));
assign g4233 = ((~g3698));
assign II12511 = ((~g7733));
assign gbuf8 = (g1956);
assign II11109 = ((~g6464));
assign II6163 = ((~g2547));
assign II5618 = ((~g1766))|((~g1771));
assign g4192 = ((~II7393));
assign II8351 = ((~g4794));
assign II10689 = ((~g6059));
assign II15229 = ((~g9968));
assign II13394 = ((~g8137));
assign g4106 = (g3284&g686);
assign g7986 = ((~g7011))|((~g6995))|((~g6984))|((~g7550));
assign g2543 = ((~II5662));
assign II15415 = ((~g10075));
assign II6388 = ((~g2329));
assign g11335 = (g11279)|(g11175);
assign g4352 = ((~II7633));
assign II15632 = ((~g10184));
assign II12369 = ((~g7189));
assign g8095 = ((~g7942));
assign g7308 = ((~II11572));
assign II12357 = ((~g7147));
assign g9773 = ((~g9474));
assign g5473 = (g4268&g3518);
assign g6193 = (g2206&g5151);
assign g4391 = ((~g3638));
assign g5900 = ((~II9531));
assign g2970 = ((~II6200))|((~II6201));
assign g6062 = ((~II9699));
assign II5612 = ((~g1280))|((~II5611));
assign g9526 = ((~g9256));
assign g4347 = ((~g3880));
assign II5296 = ((~g794))|((~II5295));
assign g3408 = ((~g3108));
assign II6065 = ((~g2226));
assign g3762 = ((~II6965));
assign g2641 = ((~g1987));
assign g7310 = ((~II11578));
assign II13959 = ((~g8451));
assign g4774 = ((~II8136));
assign II14309 = ((~g8813));
assign g6955 = ((~II11103));
assign g3071 = ((~g605))|((~g2374))|((~g2382));
assign g5544 = (g1687&g4320);
assign g6092 = (g1059&g5320);
assign g9853 = (g299&g9771);
assign g3387 = ((~II6587));
assign g10379 = ((~II15861));
assign II12372 = ((~g7137));
assign g2564 = ((~g1814));
assign II5812 = ((~g2090));
assign g8974 = (g8094&g6368&g8858);
assign g6590 = ((~g5949));
assign g8989 = ((~II14388));
assign g3632 = ((~II6799));
assign II15172 = (g9843)|(g9959)|(g9861)|(g9874);
assign g4005 = ((~II7143));
assign g3323 = ((~g2157));
assign g9576 = ((~II14713));
assign g5257 = (g691&g4755);
assign II16081 = ((~g10374))|((~II16079));
assign g7217 = (g4610&g6432);
assign II11869 = ((~g6894));
assign g4455 = ((~g3543)&(~g3419)&(~g3408));
assign g9861 = (g9738&g9579);
assign II15374 = ((~g10007));
assign II6373 = ((~g2024));
assign g2088 = ((~II4911))|((~II4912));
assign g5867 = (g3440)|(g4921);
assign g10889 = ((~II16629));
assign g11293 = (g11211)|(g10818);
assign II15879 = ((~g10359))|((~II15878));
assign II14278 = ((~g8847))|((~II14277));
assign II12180 = ((~g7263));
assign g5150 = (g1275&g4678);
assign g11502 = ((~II17525));
assign II6068 = ((~g2227));
assign II12460 = ((~g7569));
assign g7622 = ((~g7067));
assign II11778 = ((~g7210));
assign g8776 = (g5510)|(g8655);
assign g10801 = ((~II16507));
assign g5008 = (g1292&g4507);
assign g6069 = ((~II9706));
assign g11519 = (g1317&g3015&g11492);
assign II16258 = ((~g10555));
assign II16145 = (g10366&g10447&g10446);
assign II16950 = ((~g11081));
assign g6908 = (g6345)|(g4229);
assign g7301 = (g7140)|(g6327);
assign II15051 = (g7853)|(g9673)|(g9624)|(g9785);
assign g2302 = ((~g29));
assign g11466 = ((~II17435));
assign II17591 = ((~g11514));
assign g8160 = ((~II13057));
assign g10596 = ((~II16269));
assign g9150 = (g8882&g4805);
assign g6528 = (g5756)|(g4999);
assign II5840 = ((~g2432));
assign II16863 = ((~g10972));
assign g7993 = ((~II12813));
assign II8858 = ((~g4506));
assign II10412 = ((~g5821));
assign g7976 = ((~II12776));
assign g9881 = ((~g9516)&(~g9536)&(~g9573)&(~II15054));
assign g9932 = (g9911&g9624);
assign II17334 = ((~g11360));
assign g2451 = ((~g248));
assign g8020 = ((~II12862));
assign II15409 = ((~g10065));
assign II7420 = ((~g4167));
assign g6525 = (g5995&g3102);
assign g11315 = ((~II17108));
assign II15536 = ((~g10111));
assign g9847 = (g290&g9766);
assign g8048 = (g7558&g5919);
assign g7814 = ((~II12607));
assign g5005 = (g1490&g4640);
assign g2130 = ((~II5057));
assign II16537 = ((~g10721));
assign II5525 = ((~g589));
assign g11178 = (g516&g11112);
assign II13560 = ((~g722))|((~II13559));
assign g8759 = (g7437&g8677);
assign g7068 = (g5912&g6586);
assign g5082 = ((~g4840));
assign II7935 = ((~g3440));
assign g6445 = ((~II10367));
assign g10276 = ((~II15672));
assign g11302 = (g5508&g11244);
assign II13010 = ((~g8047));
assign g4437 = ((~g3345));
assign g6249 = ((~II10006));
assign g11647 = (g6622)|(g11637);
assign g6756 = (g3010&g5877);
assign g8029 = ((~II12871));
assign g6632 = (g61&g6190);
assign II13530 = ((~g704))|((~II13529));
assign g4977 = (g4567&g4807);
assign g8410 = (g713&g8143);
assign g10446 = ((~g10443))|((~g5350));
assign g11322 = ((~II17121));
assign g2642 = ((~g1988));
assign II9665 = ((~g5174));
assign g9341 = ((~II14528));
assign g6169 = ((~II9896));
assign g5626 = (g1633&g4557);
assign g2349 = ((~II5421));
assign g3627 = ((~II6784));
assign g3462 = ((~g2187)&(~g2795));
assign g8499 = (g8377&g4737);
assign g9453 = ((~g9100));
assign g7638 = (g7265)|(g6488);
assign g3426 = ((~g3121));
assign II14391 = ((~g8928));
assign g10797 = (g6206)|(g10766);
assign II13482 = ((~g8193));
assign II8396 = ((~g4255));
assign g5403 = (g4486)|(g3695);
assign g6700 = ((~g5949));
assign II12026 = ((~g7119));
assign g10655 = (g10561)|(g7389);
assign g6897 = (g6771)|(g6240);
assign g11099 = (g382&g10885);
assign g7182 = (g1878&g6720);
assign II6477 = ((~g2069));
assign g11511 = ((~II17552));
assign II9191 = ((~g5546));
assign g5944 = (g1796&g5233);
assign g10094 = ((~II15329));
assign g6237 = ((~II9984));
assign g4474 = ((~g3820));
assign II15181 = ((~g9968));
assign g7820 = (g1896&g7479);
assign g6080 = (g5249)|(g4512);
assign g4505 = (g354&g3586);
assign II6343 = ((~g1963));
assign g4345 = (g1169&g3730);
assign II13642 = ((~g8378));
assign II11515 = ((~g6589));
assign g11418 = ((~II17306))|((~II17307));
assign g5507 = (g4310&g3528);
assign g8209 = (g4094&g3792&g7980);
assign g8791 = (g8641&g8721);
assign g8271 = ((~II13185));
assign g3518 = ((~g3164));
assign II16632 = ((~g10861));
assign II9807 = ((~g5419));
assign II9443 = ((~g5557));
assign g8700 = ((~g8574));
assign II11584 = ((~g6827));
assign II5024 = ((~g995))|((~II5023));
assign II9308 = ((~g5494));
assign II12103 = ((~g6859));
assign II11794 = ((~g7188));
assign g5480 = (g4279&g3519);
assign g2041 = ((~g1791));
assign II16814 = ((~g10910));
assign g10312 = (g10220&g9094);
assign g5884 = ((~II9505));
assign II12919 = ((~g8003));
assign g2649 = ((~g2005));
assign g8334 = ((~II13382));
assign g10157 = ((~II15467));
assign g6800 = ((~II10810));
assign g6087 = (g1056&g5320);
assign g6216 = (g2232&g5151);
assign II6187 = ((~g2511))|((~II6186));
assign II10123 = ((~g5676));
assign g5423 = ((~g4300));
assign II16001 = ((~g2683))|((~II15999));
assign II11807 = ((~g6854));
assign II7726 = ((~g3378));
assign g7332 = ((~II11644));
assign II7318 = ((~g3266));
assign g11063 = ((~g10974));
assign g10267 = ((~g10130));
assign g2985 = ((~II6217));
assign g5096 = ((~g4840));
assign II7800 = ((~g3791));
assign g8964 = (g8255&g6368&g8849);
assign II13332 = ((~g8206));
assign g6036 = ((~II9647));
assign g5114 = ((~II8506));
assign g7092 = (g6540)|(g5902);
assign II12813 = ((~g7688));
assign g10284 = ((~g10167));
assign g2493 = ((~g1834))|((~g1840));
assign g11552 = (g2677&g11519);
assign g5816 = ((~II9424));
assign g9431 = ((~g9085));
assign g6917 = ((~II11029));
assign g7380 = ((~g7279));
assign II8676 = ((~g4374))|((~g1027));
assign g11635 = ((~II17719));
assign II5034 = ((~g1015))|((~g1019));
assign g3909 = ((~g2920));
assign g8585 = ((~II13828));
assign g6674 = ((~II10639));
assign g2264 = (g1771&g1766);
assign g8154 = (g7891)|(g6879);
assign g8971 = (g8081&g6764&g8858);
assign II5847 = ((~g2275));
assign II13559 = ((~g722))|((~g8263));
assign g4424 = ((~g3688));
assign g7673 = ((~II12296));
assign II11061 = ((~g6641));
assign II13283 = ((~g1927))|((~g8159));
assign g7436 = ((~g7227));
assign g4441 = ((~g3914));
assign II11916 = ((~g1494))|((~II11914));
assign g8819 = (g7957)|(g8734);
assign g6947 = ((~II11085));
assign g2120 = ((~II5035))|((~II5036));
assign g4868 = (g1027&g3914);
assign II16105 = ((~g10382));
assign g11640 = (g11613&g7900);
assign g7387 = ((~II11770));
assign g9827 = ((~II14982));
assign II12472 = ((~g7539));
assign g2846 = ((~II5970));
assign g5899 = ((~g5361));
assign II13624 = ((~g8320));
assign g7953 = ((~g7395))|((~g7390))|((~g7380))|((~g7369));
assign g2560 = ((~II5684));
assign II6812 = ((~g3290));
assign g2258 = ((~II5289));
assign g7688 = ((~g7148));
assign g2395 = ((~g231));
assign II10789 = ((~g5867));
assign g10069 = ((~II15296));
assign g10040 = ((~II15247));
assign g2346 = ((~II5414));
assign g5535 = (g4327&g3544);
assign II14672 = ((~g9261));
assign g2210 = ((~g103));
assign g6078 = (g4503)|(g5256);
assign II16507 = ((~g10712));
assign II14494 = ((~g8887));
assign g5538 = (g1669&g4313);
assign g9205 = (g6454&g8957);
assign g7594 = ((~II12120));
assign g8928 = ((~II14257));
assign II16366 = ((~g10591));
assign g3440 = ((~g3041));
assign g10459 = ((~II15968));
assign g5252 = ((~g4640));
assign g11421 = ((~II17318));
assign II5833 = ((~g2103));
assign II6001 = ((~g2548));
assign g7902 = (g7661&g6587);
assign g10531 = ((~g10471));
assign II12544 = ((~g7669));
assign g6648 = ((~II10607));
assign g7944 = ((~g7410));
assign II7707 = ((~g3370));
assign g6303 = ((~II10168));
assign II13886 = ((~g8532))|((~g1440));
assign II10858 = ((~g6688));
assign g9645 = (g1203&g9111);
assign g10542 = ((~II16193));
assign g9596 = (g2649&g9010);
assign II16938 = ((~g11086));
assign g2037 = ((~g1771));
assign g11073 = ((~g10913));
assign g8419 = ((~II13571));
assign g10335 = ((~II15787));
assign g6696 = (g5504&g5850);
assign g6575 = ((~g5949));
assign g9473 = ((~g9103));
assign g8299 = ((~II13255));
assign II7260 = ((~g2844));
assign g3060 = ((~g2135));
assign g6652 = ((~II10613));
assign g11174 = (g496&g11112);
assign g10772 = (g10655&g4840);
assign g11110 = ((~g10974));
assign g6291 = ((~II10132));
assign II9273 = ((~g5091));
assign g5587 = (g4714)|(g3904);
assign II8514 = ((~g4873))|((~II8513));
assign g1992 = ((~g782));
assign II12307 = ((~g7245));
assign II5460 = ((~g1240))|((~II5459));
assign g4444 = ((~II7800));
assign II9399 = ((~g5013));
assign g3087 = ((~II6288))|((~II6289));
assign II14537 = ((~g9308));
assign g9851 = (g296&g9770);
assign g6760 = (g786&g6221);
assign II14528 = ((~g9270));
assign II5111 = ((~g39));
assign g3997 = ((~II7131));
assign II17261 = ((~g11346));
assign g9944 = (g9924&g9392);
assign g5168 = (g1512&g4679);
assign g11340 = (g11285&g4424);
assign g7770 = ((~II12475));
assign II8180 = ((~g1786))|((~II8178));
assign g2773 = ((~II5858));
assign g6596 = ((~II10566));
assign g8568 = ((~II13797));
assign g5843 = ((~II9458));
assign g4580 = ((~g3880));
assign g8006 = ((~g5552))|((~g7717));
assign II15992 = ((~g10422))|((~g2677));
assign g8423 = ((~II13583));
assign g11349 = (g11288&g7964);
assign g2821 = ((~II5929));
assign g7790 = ((~II12535));
assign II10370 = ((~g5857));
assign g5648 = ((~II9105));
assign II15595 = ((~g10165));
assign g8752 = ((~g8635));
assign II15817 = ((~g10199));
assign g2880 = ((~II6028));
assign II13117 = ((~g7904));
assign g6855 = (g1964&g6392);
assign g9924 = (g9866)|(g9709);
assign g4269 = (g1015&g3914);
assign II4985 = ((~g999))|((~g1003));
assign g7130 = (g6041&g6697);
assign II9290 = ((~g5052));
assign g2760 = (g981&g2091);
assign g4177 = ((~II7348));
assign g10892 = ((~II16638));
assign II6395 = ((~g2334));
assign II10592 = ((~g5865));
assign g11556 = (g2701&g11519);
assign g10343 = ((~II15795));
assign II12424 = ((~g7635));
assign g2755 = ((~II5833));
assign II8771 = ((~g4619))|((~II8770));
assign II15704 = ((~g10238));
assign g5721 = (g1577&g5143);
assign g2862 = ((~g2315)&(~g2305));
assign g7476 = ((~g6933));
assign g5597 = ((~II9023));
assign g4389 = (g3529&g3092);
assign II14687 = ((~g9258));
assign g4748 = ((~g3546));
assign II14473 = ((~g8921));
assign II15176 = (g8176)|(g9910)|(g9897)|(g9836);
assign g4735 = ((~g3546));
assign g4078 = ((~II7205));
assign g4280 = ((~g4013));
assign g3351 = ((~II6535));
assign II13666 = ((~g8292));
assign II6917 = ((~g2832));
assign g6881 = ((~II10971));
assign II4978 = ((~g411))|((~g333));
assign g10382 = ((~g10314)&(~g2998));
assign g3378 = ((~II6572));
assign g5615 = ((~II9043));
assign g2103 = ((~II4961));
assign g11619 = ((~II17675));
assign II13030 = ((~g8052));
assign II4971 = ((~g991))|((~g995));
assign g7736 = (g6951&g3880);
assign g11083 = ((~g10913));
assign g4439 = ((~II7793));
assign g7479 = ((~II11873));
assign g11652 = ((~II17758));
assign g3636 = ((~II6815));
assign II14179 = ((~g8785));
assign g5590 = (g4718)|(g4723);
assign g2732 = ((~II5792));
assign g8614 = (g8365)|(g8510);
assign g8178 = ((~II13083));
assign II11505 = ((~g6585));
assign g11043 = ((~II16790));
assign g4290 = ((~g3586));
assign g8352 = ((~II13436));
assign g10199 = ((~g10172));
assign g4791 = ((~II8161));
assign g2251 = ((~g731));
assign g5827 = ((~II9443));
assign g6387 = ((~g6121));
assign II6690 = ((~g2743));
assign g7990 = ((~g7011))|((~g6995))|((~g7562))|((~g7550));
assign II10898 = ((~g6735));
assign g2076 = ((~II4886));
assign g7799 = ((~II12562));
assign g10497 = (g5052)|(g10396);
assign g9601 = (g922&g9192);
assign g5877 = (g4921&g639);
assign II6907 = ((~g2994));
assign g3380 = ((~II6576));
assign g7765 = ((~II12460));
assign g3306 = ((~II6477));
assign II9905 = ((~g5300));
assign II7429 = ((~g3344));
assign II15517 = ((~g10051));
assign g6452 = ((~II10384));
assign g8706 = (g7602&g8589);
assign g6410 = (g2804&g5759);
assign g9967 = (g9957&g9536);
assign g5353 = ((~II8820));
assign g10705 = (g10564&g4840);
assign II9652 = ((~g5426));
assign g8424 = ((~II13586));
assign g8432 = (g8389)|(g8072);
assign g10538 = ((~II16181));
assign II16941 = ((~g11076));
assign g8732 = (g8624&g7919);
assign g2163 = ((~II5092));
assign g2808 = ((~g2156));
assign g6095 = (g1062&g5320);
assign g4996 = (g1428&g4682);
assign II14376 = ((~g8959));
assign g7844 = ((~II12631));
assign g7703 = ((~g7085));
assign g11035 = ((~II16766));
assign II15589 = ((~g10161));
assign g6661 = (g73&g6219);
assign g6267 = ((~II10060));
assign g7582 = ((~II12061))|((~II12062));
assign g4099 = (g770&g3281);
assign g8480 = ((~II13682));
assign g5284 = ((~g4376));
assign II10189 = ((~g6112));
assign g4673 = ((~g4013));
assign II6538 = ((~g2827));
assign g2502 = ((~II5579));
assign II11668 = ((~g7043));
assign II5136 = ((~g521))|((~II5135));
assign g4142 = ((~II7288));
assign II11909 = ((~g1474))|((~II11907));
assign II11671 = ((~g7047));
assign g5790 = ((~II9388));
assign g5180 = (g4541&g4533);
assign II13732 = ((~g8291));
assign II10946 = ((~g6548));
assign II12822 = ((~g7677));
assign II7465 = ((~g3726));
assign II9150 = ((~g5012));
assign g4125 = ((~II7272));
assign II13506 = ((~g8247))|((~II13504));
assign II11650 = ((~g6938));
assign g10035 = ((~II15241));
assign g2305 = (II5351)|(II5352);
assign g10131 = ((~II15395));
assign II5795 = ((~g2462));
assign g4885 = ((~II8228));
assign II5713 = ((~g2436));
assign g5187 = ((~II8590))|((~II8591));
assign II12993 = ((~g8044));
assign g5784 = ((~II9380));
assign g9358 = (g1318&g9151);
assign g8220 = ((~g7826));
assign g11159 = ((~g10950));
assign g7530 = ((~II11926));
assign II5570 = (g416)|(g411)|(g406)|(g401);
assign g7964 = ((~g7651));
assign g10511 = ((~g10438))|((~g6032));
assign g7995 = ((~II12817));
assign g5730 = ((~II9282));
assign g8386 = (g6085&g8219);
assign II13678 = ((~g8306));
assign g4367 = ((~II7662));
assign II9188 = ((~g4908));
assign g9588 = (g3272&g9173);
assign g8120 = (g1909&g7944);
assign g11618 = ((~II17672));
assign g2217 = ((~II5192));
assign g8347 = ((~II13421));
assign g6353 = (g299&g5895);
assign g6735 = ((~II10736));
assign g7981 = ((~g7624));
assign g6983 = (g6592&g3105);
assign II4910 = ((~g386))|((~g318));
assign II16479 = ((~g10767));
assign II16595 = ((~g10783));
assign II15427 = ((~g10088));
assign II11166 = ((~g6480));
assign g7524 = ((~II11915))|((~II11916));
assign II8973 = ((~g4488));
assign g2947 = ((~II6137))|((~II6138));
assign II8642 = ((~g516))|((~II8640));
assign g11504 = ((~II17531));
assign II7017 = ((~g3068));
assign g8155 = ((~II13048));
assign g7504 = (g7148&g2847);
assign g4241 = ((~g3664));
assign g5862 = ((~II9479));
assign II8577 = ((~g496))|((~II8575));
assign g2201 = ((~g102));
assign g9694 = (g278&g9432);
assign g7187 = ((~II11405));
assign g10323 = ((~II15763));
assign g6120 = ((~II9813));
assign gbuf1 = (g883);
assign II4786 = ((~g109));
assign g8269 = (g7892)|(g3429);
assign g8547 = (g8307&g7693);
assign II6671 = ((~g2757));
assign g11235 = (g5443&g11107);
assign g9258 = ((~g8892));
assign g10672 = (g10579&g9449);
assign g7851 = ((~g7479));
assign g4313 = ((~g3586));
assign g7445 = ((~II11845));
assign II5998 = ((~g2197));
assign g4963 = ((~II8337));
assign II15744 = ((~g10261));
assign g2055 = ((~g1950));
assign g2952 = ((~g2455));
assign g5795 = (g1543&g5251);
assign g10690 = (g10616&g3863);
assign g7034 = ((~II11191));
assign g9010 = (g6454&g8930);
assign II15717 = ((~g10231))|((~II15716));
assign II12150 = ((~g7074));
assign II9598 = ((~g5120));
assign g3766 = ((~g2439))|((~g3222))|((~g2493));
assign g11439 = ((~II17368));
assign g5701 = ((~II9240));
assign g8135 = (g1945&g7956);
assign g5484 = (g1896&g4256);
assign g11399 = ((~II17240));
assign g3937 = ((~II7086));
assign g8169 = (g5265&g7853);
assign II6367 = ((~g2045));
assign g11337 = (g11282)|(g11177);
assign g10236 = ((~g10190));
assign g4711 = ((~II8061));
assign g2436 = ((~II5525));
assign g1991 = ((~g778));
assign II13255 = ((~g8270));
assign g8739 = ((~g8640));
assign g5270 = ((~g4367));
assign g8888 = ((~II14232));
assign g3103 = ((~g2391));
assign g7273 = ((~g6365));
assign g9917 = (g9856)|(g9695);
assign II6738 = ((~g3113));
assign II4820 = ((~g865));
assign g4105 = ((~II7249));
assign II14055 = ((~g8650));
assign g9993 = ((~II15193));
assign g3226 = ((~II6403));
assign g10256 = ((~g10140));
assign II13941 = ((~g8488));
assign g7225 = (g6666)|(g6079);
assign g4449 = ((~g4144));
assign g11227 = (g11151)|(g11010);
assign g4775 = ((~II8139));
assign g3110 = ((~g2482));
assign g5770 = (g4466&g5128);
assign II12496 = ((~g7724));
assign II10541 = ((~g6176));
assign g2240 = ((~g88));
assign II4964 = ((~g406))|((~g330));
assign g5300 = ((~II8771))|((~II8772));
assign II16217 = ((~g10501));
assign g7545 = ((~II11967));
assign g6149 = ((~II9866));
assign II12174 = ((~g6939));
assign II12053 = ((~g6928));
assign II5325 = ((~g1341))|((~II5323));
assign g8311 = ((~II13317));
assign g7134 = (g5587&g6354);
assign g7291 = (g7050)|(g6317);
assign II6077 = ((~g2349));
assign II7677 = ((~g3735));
assign g9723 = (g9620)|(g9652)|(g9391)|(II14858);
assign II17305 = ((~g11381))|((~g11377));
assign II8164 = ((~g3566));
assign g10228 = ((~II15604));
assign II7564 = ((~g654))|((~II7562));
assign g11577 = ((~II17613));
assign II13837 = ((~g8488));
assign g7558 = ((~II12003))|((~II12004));
assign II10293 = ((~g5863));
assign g10766 = (g10646&g4840);
assign II6733 = ((~g3321));
assign g7758 = ((~II12439));
assign g8463 = (g8301&g7410);
assign II5224 = ((~g61));
assign II17104 = ((~g11223));
assign g6273 = ((~II10078));
assign g6814 = ((~II10852));
assign g2639 = ((~II5754));
assign II7223 = ((~g2981))|((~g1781));
assign II17249 = ((~g11342));
assign g5739 = (g1607&g5185);
assign g8948 = ((~II14299));
assign II13992 = ((~g8688))|((~II13990));
assign II16038 = ((~g10427))|((~II16037));
assign II10885 = ((~g6332));
assign g11026 = (g386&g10974);
assign II11543 = ((~g6881));
assign II14452 = ((~g8922));
assign g7557 = ((~II11996))|((~II11997));
assign II14123 = ((~g8767));
assign g5919 = (g5216&g2965);
assign g2748 = ((~II5812));
assign g4296 = ((~II7559));
assign II11152 = ((~g6469));
assign g10243 = ((~II15635));
assign g10492 = ((~II16111));
assign g4231 = (g3991)|(g3998);
assign g6339 = ((~II10240));
assign g8571 = ((~II13806));
assign II14083 = ((~g8747));
assign g5941 = ((~II9571));
assign g10315 = ((~g10243));
assign g11561 = (g11518&g3015);
assign II7875 = ((~g4109))|((~g810));
assign g3222 = ((~g2557))|((~g1814))|((~g1834));
assign g8464 = (g8302&g7416);
assign g10674 = ((~g10584));
assign g6278 = ((~II10093));
assign g5666 = ((~II9159));
assign II10589 = ((~g5763));
assign II16289 = ((~g10541));
assign II15219 = (g8172)|(g9907)|(g9936)|(g9833);
assign II13236 = ((~g8245));
assign g4781 = ((~II8147));
assign g6103 = ((~II9766));
assign II16461 = ((~g10735));
assign II5002 = ((~g1173));
assign II11973 = ((~g7001))|((~g1462));
assign g9532 = ((~II14681));
assign g6343 = ((~II10248));
assign g4331 = ((~II7606));
assign g7660 = (g7059)|(g6583);
assign II9946 = ((~g5233))|((~g1796));
assign II6443 = ((~g2363));
assign g4214 = ((~II7459));
assign g2963 = ((~II6187))|((~II6188));
assign g2828 = ((~II5940));
assign g8263 = (g8032)|(g7720);
assign g4167 = ((~II7318));
assign gbuf6 = (g113);
assign g10936 = (g5170)|(g10808);
assign g3976 = ((~II7109));
assign g6054 = (g5199)|(g4483);
assign g9615 = ((~g9052)&(~g9030));
assign g4279 = ((~II7536));
assign II15441 = ((~g10035))|((~g10122));
assign g6001 = ((~II9625));
assign g10200 = ((~g10169));
assign g10248 = ((~g10134));
assign g3695 = (g1712&g3015);
assign g10852 = ((~g10740));
assign g8145 = ((~II13030));
assign II13242 = ((~g8267));
assign g2778 = ((~g2276));
assign g8939 = (g8791)|(g8701);
assign g6874 = ((~II10958));
assign g2194 = ((~g47));
assign g4458 = ((~II7817));
assign g6254 = ((~II10021));
assign II16468 = ((~g10716))|((~II16467));
assign g11587 = (g1327&g11546);
assign II4920 = ((~g260));
assign g4726 = ((~g3546));
assign II4935 = ((~g585));
assign II5878 = ((~g2120))|((~g2115));
assign II9135 = ((~g5198));
assign g10484 = (g9317)|(g10400);
assign g9490 = ((~g9324));
assign g8125 = ((~II12986));
assign g10128 = ((~II15386));
assign g7103 = ((~II11338));
assign g10874 = ((~II16592));
assign g7617 = ((~II12199));
assign g2801 = ((~g2117));
assign g10665 = ((~II16331))|((~II16332));
assign g6540 = (g1223&g6072);
assign g6570 = ((~g5949));
assign g9941 = (g9921&g9367);
assign g3370 = ((~II6560));
assign g2604 = ((~II5713));
assign g10733 = (g5227)|(g10674);
assign II9415 = ((~g5047));
assign g10759 = (g10698&g10697);
assign g8104 = (g6218&g7880);
assign g7413 = ((~g7197));
assign g4083 = ((~II7216));
assign g9292 = (g8878&g5708);
assign g2173 = ((~II5120));
assign II10553 = ((~g6192));
assign II10891 = ((~g6334));
assign g11473 = ((~II17456));
assign g4876 = (g1086&g3638);
assign II5478 = ((~g1212));
assign g6071 = (g5228)|(g4505);
assign II15787 = ((~g10269));
assign II12601 = ((~g7629));
assign g3863 = (g3323&g2728);
assign g8409 = ((~II13530))|((~II13531));
assign g3039 = ((~g2310));
assign g9815 = ((~g9392)&(~g9367));
assign g4497 = (g351&g3586);
assign g5089 = ((~g4840));
assign g5109 = ((~II8495));
assign g2353 = (g1403)|(g1407)|(g1411)|(g1415);
assign II11617 = ((~g6839));
assign g7375 = (g7230)|(g6745);
assign g5104 = (g1796&g4608);
assign g11447 = ((~II17390));
assign g11205 = ((~g11112));
assign g4807 = (g3015&g1289&g3937);
assign g7748 = ((~II12409));
assign g5425 = ((~g4300));
assign g7406 = ((~II11786));
assign g3485 = ((~g2662));
assign g4323 = ((~g4130));
assign II15983 = ((~g10414));
assign II11572 = ((~g6822));
assign g5633 = ((~g4388));
assign g9103 = ((~g8892));
assign II9833 = ((~g5197));
assign g8473 = ((~II13669));
assign II8678 = ((~g1027))|((~II8676));
assign II7710 = ((~g3749));
assign g10292 = ((~II15698));
assign II8268 = ((~g4674));
assign g2965 = ((~II6196));
assign g2873 = ((~II6019));
assign g8871 = ((~II14185));
assign g10934 = ((~g10827));
assign II6138 = ((~g378))|((~II6136));
assign II13188 = ((~g8171));
assign g4318 = ((~g4130));
assign g6836 = ((~II10888));
assign g4007 = (g2683&g2276);
assign II7513 = ((~g4144));
assign g6667 = ((~II10630));
assign II12878 = ((~g7638));
assign g7325 = ((~II11623));
assign II11146 = ((~g6439));
assign g7004 = ((~II11143));
assign g10299 = (g8892&g10217);
assign II7210 = ((~g2798));
assign g7924 = ((~g7470));
assign II13909 = ((~g1432))|((~II13907));
assign g11253 = (g981&g11072);
assign II7363 = ((~g4005));
assign g4376 = ((~II7691));
assign g8251 = ((~II13166));
assign g5853 = (g5044&g1927);
assign II9123 = ((~g4890));
assign g2070 = ((~g213));
assign g6164 = ((~g5426));
assign II10156 = ((~g6100));
assign II7732 = ((~g3758));
assign g11023 = (g440&g10974);
assign g2081 = (g932&g928);
assign g8435 = (g8403)|(g8075);
assign g10862 = (g5524)|(g10746);
assign II6424 = ((~g2462));
assign g4767 = ((~II8123));
assign g3318 = ((~g2245));
assign g10513 = ((~g10441))|((~g5345));
assign g6552 = ((~g5733));
assign g10820 = ((~II16528));
assign g11223 = (g11147)|(g11008);
assign II17447 = ((~g11457));
assign g9079 = ((~g8892));
assign g7922 = ((~II12712));
assign g1962 = ((~g27));
assign II12930 = ((~g7896));
assign II7757 = ((~g3767));
assign II10804 = ((~g6388));
assign II13307 = ((~g8190))|((~g617));
assign g5573 = ((~g4117)&(~g4432));
assign g11623 = ((~II17687));
assign II14519 = ((~g9106));
assign g8816 = (g7951)|(g8731);
assign g5619 = ((~g4840));
assign g10202 = ((~g10171));
assign II7462 = ((~g3721));
assign g6245 = (g575&g5098);
assign g4562 = ((~II7973));
assign II17438 = ((~g11444));
assign II6799 = ((~g2750));
assign g8743 = ((~g8617))|((~g6971))|((~g6964));
assign g8320 = ((~II13344));
assign g10422 = ((~g10289)&(~g4620));
assign g9778 = ((~g9474));
assign g6702 = ((~g5949));
assign II12265 = ((~g7211));
assign II14130 = ((~g8769));
assign II12439 = ((~g7663));
assign g3205 = ((~g1814))|((~g2571));
assign g6934 = (g6363)|(g5720);
assign g4253 = (g1074&g3638);
assign II8885 = ((~g4548));
assign II11981 = ((~g6957))|((~II11980));
assign g2299 = ((~g1707));
assign II6771 = ((~g3257))|((~II6770));
assign g10429 = ((~g10326)&(~g3507));
assign II7387 = ((~g4083));
assign g3413 = ((~g2896));
assign g10728 = (g4973)|(g10642);
assign g4201 = ((~II7420));
assign g11395 = ((~II17228));
assign g7258 = (g6549)|(g5913);
assign g4535 = ((~g3946));
assign g8825 = ((~g8502))|((~g8738))|((~g8506));
assign II10192 = ((~g6115));
assign g5802 = (g5601)|(g4837);
assign g7421 = ((~II11807));
assign II5886 = (g174&g170&g2249&g2254);
assign g2960 = ((~II6173));
assign g9959 = (g9950&g9536);
assign II17384 = ((~g11437));
assign II12532 = ((~g7594));
assign g9522 = (g9173)|(g9125);
assign g4088 = ((~II7224))|((~II7225));
assign g9528 = (g9151)|(g9125)|(g9111);
assign g8955 = (g8110&g6368&g8828);
assign II9612 = ((~g5149));
assign g4518 = (g452&g3975);
assign g9411 = (g1724&g9052);
assign g7717 = ((~g6863))|((~g3206));
assign II11623 = ((~g6841));
assign g7612 = ((~II12186));
assign g8474 = (g8383&g5285);
assign g2655 = ((~g2013));
assign g10487 = ((~II16098));
assign II14585 = (g8995)|(g9205)|(g9192);
assign g9899 = (g9889&g9367);
assign II5265 = ((~g461))|((~II5263));
assign II16178 = ((~g10490));
assign g8182 = ((~II13099));
assign g2794 = (II5886&II5887);
assign g6256 = ((~II10027));
assign g2236 = ((~II5230))|((~II5231));
assign g4209 = ((~II7444));
assign g5688 = ((~II9213));
assign g9854 = (g9730&g9566);
assign g3331 = ((~II6510));
assign g7127 = (g6663&g2241);
assign g10390 = ((~g10309));
assign II13561 = ((~g8263))|((~II13559));
assign g10143 = ((~II15427));
assign II8116 = ((~g3627));
assign g7123 = ((~II11360));
assign g10707 = (g5545)|(g10686);
assign g4721 = ((~g3546));
assign g11165 = (g476&g11112);
assign g5645 = ((~II9096));
assign II15278 = ((~g10033));
assign II6616 = ((~g3186));
assign g9671 = ((~II14802));
assign g7720 = (g727&g7232);
assign II11211 = ((~g6527));
assign II8989 = ((~g4746));
assign g5043 = ((~g4840));
assign g3730 = ((~g3015));
assign g11608 = (g11587)|(g11558);
assign g8482 = ((~g8329));
assign II10437 = ((~g5755));
assign g11258 = (g11235)|(g11020);
assign g6718 = ((~g5949));
assign g2225 = ((~II5210));
assign II14793 = ((~g9269));
assign g4052 = (g2862)|(g2515);
assign g4073 = (g3200&g3222);
assign g2180 = ((~II5136))|((~II5137));
assign II11338 = ((~g6680));
assign II14109 = ((~g8765));
assign g6537 = (g5781)|(g5005);
assign g4011 = ((~II7151));
assign g7788 = ((~II12529));
assign II5593 = ((~g1703))|((~II5591));
assign g7738 = (g7200)|(g6738);
assign g11548 = ((~g11519));
assign II16644 = ((~g10865));
assign g5123 = (g1618&g4669);
assign g8079 = ((~II12939));
assign II11956 = ((~g6912));
assign II9699 = ((~g5426));
assign g5789 = (g1561&g5232);
assign g6517 = ((~II10434));
assign g10608 = ((~II16283));
assign g2765 = ((~g2184));
assign g9553 = ((~II14694));
assign g6325 = (g1245&g5949);
assign II7236 = ((~g3219));
assign g6046 = ((~II9669));
assign g10271 = ((~II15665));
assign g8771 = (g5483)|(g8652);
assign g8617 = ((~g8465));
assign II13803 = ((~g8476));
assign II11005 = ((~g6386));
assign g8008 = ((~II12846));
assign g5419 = ((~II8858));
assign g6423 = (g4348&g5784);
assign g9353 = ((~II14564));
assign g10680 = (g10564&g3586);
assign g5902 = (g2555&g4977);
assign g11318 = (g11228)|(g11104);
assign II15448 = ((~g10056));
assign II5854 = ((~g2523));
assign g7705 = (g6853&g4328);
assign II14805 = ((~g9360));
assign II14385 = ((~g8890));
assign II12274 = ((~g7110));
assign II14955 = ((~g9765));
assign II6921 = ((~g2839));
assign g4368 = ((~II7665));
assign g6113 = ((~II9792));
assign II10535 = ((~g5867));
assign II12165 = ((~g6882));
assign II7339 = ((~g4004));
assign II14209 = ((~g8824))|((~g599));
assign g5126 = (g3076&g4638);
assign II11447 = ((~g6431));
assign g2094 = ((~II4924));
assign II16255 = ((~g10554));
assign II13900 = ((~g8520))|((~g1428));
assign g7880 = ((~g7479));
assign g4891 = (g631&g4739);
assign g11622 = ((~II17684));
assign g8601 = ((~g8477));
assign gbuf13 = (g1217);
assign g2186 = ((~g90));
assign g4325 = (g1166&g3682);
assign II12514 = ((~g7735));
assign g5691 = ((~g5236));
assign II9311 = ((~g4915));
assign g5896 = ((~II9525));
assign II13068 = ((~g7906));
assign g7340 = ((~II11668));
assign g5674 = (g148&g5361);
assign II8545 = ((~g486))|((~II8543));
assign g7366 = ((~II11746));
assign II10477 = ((~g6049));
assign II12113 = ((~g7093))|((~g162));
assign g7220 = ((~II11456));
assign g5679 = ((~II9194));
assign II8487 = ((~g4526));
assign g6711 = ((~g5949));
assign g10552 = ((~II16217));
assign g7059 = (g6078&g6714);
assign g6470 = (g5699)|(g4960);
assign g5236 = ((~g4361));
assign g4484 = (g1137&g3909);
assign g7322 = ((~II11614));
assign g2232 = ((~II5221));
assign II10710 = ((~g6088));
assign g3263 = (g2503&g2328);
assign g7204 = (g6645)|(g6062);
assign g2998 = ((~g2462));
assign g7271 = (g5028&g6499);
assign g1984 = ((~g758));
assign g5176 = ((~g4682));
assign g7727 = ((~II12366));
assign II16052 = ((~g837))|((~II16051));
assign II5620 = ((~g1771))|((~II5618));
assign g11481 = (g6624)|(g11458);
assign g7319 = ((~II11605));
assign g4261 = (g1019&g3914);
assign g8608 = ((~g8482));
assign g7031 = ((~g6413));
assign g10435 = ((~g10332)&(~g3507));
assign II15559 = ((~g10094));
assign II9571 = ((~g5509));
assign g4243 = ((~g3524));
assign g4618 = ((~g3829));
assign II12261 = ((~g7078));
assign II15431 = ((~g10047))|((~II15430));
assign g4198 = ((~II7411));
assign II5818 = ((~g2098));
assign g2433 = ((~II5517))|((~II5518));
assign g10716 = (g10497&g10675);
assign II7776 = ((~g3773));
assign II6988 = ((~g2760))|((~g986));
assign II8211 = ((~g3566));
assign g5658 = ((~II9135));
assign II15520 = ((~g10035));
assign II17684 = ((~g11609));
assign g11478 = (g6532)|(g11455);
assign g11157 = ((~g10950));
assign g10303 = (g10208&g9076);
assign g11468 = ((~II17441));
assign II15383 = ((~g10107));
assign g8625 = ((~g8487));
assign g4903 = (g1849&g4243);
assign II9813 = ((~g5241));
assign II10971 = ((~g6344));
assign g3764 = ((~II6971));
assign g5997 = ((~II9617));
assign g9711 = (g9660)|(g9390)|(g9359)|(g9589);
assign II12454 = ((~g7544));
assign II13659 = ((~g1945))|((~g8322));
assign g10803 = ((~g10708));
assign g9656 = ((~g9010)&(~g9240)&(~g9223)&(~II14779));
assign g7900 = ((~g7712));
assign g7040 = ((~II11207));
assign g5073 = ((~g4840));
assign II11351 = ((~g6698));
assign g7805 = ((~II12580));
assign g9663 = (g959&g9223);
assign g10443 = ((~g10353)&(~g3566));
assign g10904 = ((~II16664));
assign g2837 = ((~g2130));
assign II9111 = ((~g5596));
assign g8769 = (g8629&g5151);
assign g5753 = ((~II9329));
assign g6026 = (g5507)|(g3970);
assign g8100 = ((~g7947));
assign II17353 = ((~g11381));
assign g2789 = ((~g2276));
assign II15287 = ((~g9980));
assign II9205 = ((~g5309));
assign g9563 = (g9052)|(g9030);
assign II11322 = ((~g6652));
assign II6990 = ((~g986))|((~II6988));
assign g3015 = (g2028&g2191);
assign II11360 = ((~g6351));
assign g3255 = ((~II6421));
assign II13537 = ((~g658))|((~g8157));
assign g7946 = ((~g7416));
assign II14116 = ((~g8766));
assign g6547 = ((~g5893));
assign g6235 = (g569&g5089);
assign g3819 = (g3275)|(g9);
assign II12232 = ((~g7072));
assign g9771 = ((~g9432));
assign g9757 = ((~g9454)&(~g9274)&(~g9292));
assign g4728 = ((~II8080));
assign g2480 = ((~II5561));
assign II8290 = ((~g4778));
assign g9761 = ((~g9454));
assign II10066 = ((~g5778));
assign g6060 = ((~II9695));
assign g6990 = ((~II11132));
assign g7463 = ((~g6921));
assign g9990 = ((~II15190));
assign II10456 = ((~g5844));
assign II13888 = ((~g1440))|((~II13886));
assign g8200 = (g7535)|(g8008);
assign g9731 = (g9641)|(g9364)|(g9387);
assign g10360 = ((~g10277)&(~g3566));
assign g4121 = ((~II7264));
assign g10622 = (g10543&g4525);
assign g10600 = ((~II16277));
assign g7933 = (g2814&g7450);
assign g5469 = ((~II8880));
assign g8961 = ((~II14330));
assign II5866 = ((~g2107))|((~II5865));
assign g4969 = (g1642&g4463);
assign g6502 = (g5981&g3095);
assign g8190 = ((~g6027))|((~g7978));
assign g8733 = (g8625&g7920);
assign II17271 = ((~g11388));
assign g7629 = ((~II12229));
assign g5275 = ((~g4371));
assign g8099 = ((~g7990));
assign g4495 = ((~II7886));
assign II10907 = ((~g6705));
assign g4359 = ((~g3880));
assign g5542 = ((~II8967));
assign g5720 = (g170&g5361);
assign g8546 = ((~g3983))|((~g8390));
assign g4235 = (g1011&g3914);
assign g6194 = (g554&g5043);
assign g11457 = ((~II17424));
assign g8553 = (g8405&g8015);
assign g11242 = ((~g11112));
assign g2910 = (g2424&g1660);
assign g7355 = ((~II11713));
assign II15473 = ((~g10087));
assign g9256 = (g6689&g8963);
assign g9960 = (g9951&g9536);
assign II11824 = ((~g7246));
assign II11528 = ((~g6796));
assign g10187 = ((~II15539));
assign g3536 = (g2390&g3103);
assign II15485 = ((~g10092));
assign g11146 = (g318&g10928);
assign II7956 = ((~g3428));
assign g5254 = (g4335&g4165);
assign II11464 = ((~g6443));
assign g8886 = ((~II14228));
assign g2110 = ((~II5002));
assign II12953 = ((~g8024));
assign g7590 = (g7102&g5425);
assign g10411 = (g10299)|(g9529);
assign g5471 = ((~g4370));
assign g8218 = ((~g7826));
assign II8900 = ((~g4560));
assign g8050 = (g7596&g5919);
assign II8250 = ((~g4589));
assign g9265 = ((~g8892));
assign g8987 = ((~II14382));
assign g2529 = ((~II5638));
assign g6950 = ((~II11094));
assign g5401 = ((~II8839));
assign g6067 = (g1047&g5320);
assign II12092 = ((~g6944))|((~g1490));
assign g7978 = ((~g7697))|((~g3038));
assign g3634 = ((~II6806))|((~II6807));
assign II16650 = ((~g10776));
assign g10352 = ((~II15820));
assign II6126 = ((~g1419))|((~II6124));
assign II5372 = ((~g971))|((~II5371));
assign II5210 = ((~g58));
assign g11307 = ((~II17092));
assign g10901 = ((~g10802));
assign II14555 = ((~g9009));
assign II12293 = ((~g7116));
assign g3428 = ((~II6639));
assign g7624 = ((~II12215))|((~II12216));
assign g10389 = ((~g10307));
assign g11053 = ((~g10950));
assign g10780 = (g10723&g5124);
assign II12074 = ((~g7098))|((~g174));
assign g6626 = (g5934)|(g123);
assign g7812 = ((~II12601));
assign II8527 = ((~g4879))|((~g481));
assign g5555 = (g4389)|(g4397);
assign g9938 = (g9917&g9367);
assign g11498 = ((~II17513));
assign II14910 = ((~g9532));
assign II9388 = ((~g5576));
assign II6016 = ((~g2201));
assign II5584 = ((~g1200));
assign g2245 = ((~II5254));
assign II13592 = ((~g8362));
assign g9930 = ((~II15127));
assign g9768 = ((~g9432));
assign g10047 = ((~II15266));
assign g9507 = ((~g9268));
assign II8520 = ((~g4338));
assign g6943 = ((~II11079));
assign II6630 = (g2677&g2683&g2689&g2701);
assign II4780 = ((~g872));
assign g7025 = ((~g6400));
assign g6586 = ((~g5949));
assign II5142 = ((~g639));
assign g9425 = (g1753&g9030);
assign g7106 = (g6554)|(g5917);
assign II16626 = ((~g10859));
assign II12099 = ((~g7258));
assign g8039 = (g7587&g5128);
assign g4753 = (g481&g3386);
assign g8229 = ((~g7826));
assign g11218 = (g959&g11053);
assign II6224 = ((~g2544))|((~g1346));
assign g6090 = (g553&g5627);
assign II15864 = ((~g10339));
assign II17371 = ((~g11410));
assign II9792 = ((~g5403));
assign II5765 = ((~g2004));
assign II10093 = ((~g5779));
assign g7605 = ((~II12165));
assign II11252 = ((~g6542));
assign g7822 = (g1914&g7479);
assign g4952 = (g1648&g4457);
assign II16772 = ((~g10887));
assign g7416 = ((~II11800));
assign g3621 = ((~II6754));
assign g4361 = ((~II7648));
assign II10648 = ((~g6030));
assign g2885 = ((~II6043));
assign g7209 = (g3804&g6425);
assign g8193 = (g5145)|(g7937);
assign g7350 = ((~II11698));
assign g10387 = ((~g10357));
assign II13191 = ((~g8132));
assign g10185 = ((~g10040));
assign g11426 = ((~II17331));
assign g2381 = ((~g1368));
assign II15965 = ((~g10405));
assign II10033 = ((~g5693));
assign g4300 = (g3546)|(g2391);
assign g6220 = ((~g5446));
assign II6557 = ((~g3086));
assign g5718 = ((~II9256));
assign II10904 = ((~g6558));
assign II15698 = ((~g10235));
assign II9320 = ((~g5013));
assign II10724 = ((~g6096));
assign g8115 = ((~g7953));
assign g8360 = ((~II13460));
assign g4770 = (g416&g3415);
assign II8036 = ((~g3820));
assign g7074 = ((~II11299));
assign g10774 = ((~II16458));
assign g5420 = ((~g4300));
assign g3345 = ((~II6531));
assign g10687 = ((~II16356));
assign g5349 = (g2126&g4617);
assign II11345 = ((~g6692));
assign g6479 = (g5707)|(g4968);
assign g11450 = ((~II17407));
assign g6509 = ((~II10427));
assign II5966 = ((~g2541));
assign g2101 = ((~II4951));
assign g5727 = ((~II9273));
assign II6932 = ((~g2850));
assign II17755 = ((~g11646));
assign g5470 = (g1044&g4222);
assign g7516 = ((~g7148));
assign g10577 = ((~g10526));
assign II8429 = ((~g4458));
assign g7760 = ((~II12445));
assign g4943 = ((~II8311));
assign g4587 = ((~g3829));
assign II12595 = ((~g7706));
assign g9260 = ((~g8892));
assign II12875 = ((~g7638));
assign g10795 = (g6199)|(g10764);
assign g6922 = (g6352)|(g5694);
assign g11580 = (g11413)|(g11544);
assign g5494 = ((~g4412));
assign g5215 = (g4276&g3400);
assign g8725 = ((~g8589));
assign g6284 = ((~II10111));
assign g7028 = ((~g6407));
assign II15568 = ((~g10094));
assign g6805 = ((~II10825));
assign g9884 = ((~II15063));
assign II12183 = ((~g7007));
assign g2522 = (g833)|(g829)|(II5629);
assign g7774 = ((~II12487));
assign g9702 = (g9365)|(g9647)|(II14831);
assign g8070 = (g682&g7826);
assign II14224 = ((~g8794));
assign II17191 = ((~g11315));
assign g5756 = (g1531&g5202);
assign g2396 = ((~g1389));
assign II11261 = ((~g6775))|((~g826));
assign g7061 = (g790&g6760);
assign g8404 = (g686&g8129);
assign g6320 = (g1292&g5949);
assign g9729 = (g9618)|(g9357)|(g9656);
assign g4620 = ((~II8031));
assign II10057 = ((~g5741));
assign g9097 = ((~g8892));
assign II13212 = ((~g8195));
assign g7889 = (g7615&g3814);
assign g10150 = ((~II15448));
assign II8778 = ((~g4630))|((~g1137));
assign g6404 = (g2132&g5748);
assign g10282 = ((~g10164));
assign g10119 = ((~II15365));
assign g7196 = ((~II11420));
assign g8841 = (g8605&g8704);
assign II9510 = ((~g5421));
assign g8848 = (g8715&g8713);
assign g11276 = ((~II17052))|((~II17053));
assign g4986 = (g1411&g4682);
assign g8684 = ((~II13969));
assign g10580 = ((~g10530));
assign g8062 = ((~II12904));
assign II12039 = ((~g6990))|((~II12038));
assign g10034 = ((~II15238));
assign g9511 = (g9151)|(g9125)|(g9111);
assign g7278 = ((~II11524));
assign g3394 = ((~II6598));
assign g7907 = ((~g7664));
assign g8991 = ((~II14394));
assign g4398 = ((~g3914));
assign g3810 = ((~g3228));
assign g2074 = ((~g1377));
assign II14295 = ((~g8806));
assign g11596 = ((~g11580));
assign g6929 = (g6360)|(g5704);
assign g11313 = ((~II17104));
assign g11554 = (g2689&g11519);
assign g6202 = ((~g5426));
assign g4199 = ((~II7414));
assign II6517 = ((~g3271));
assign g4182 = ((~II7363));
assign II15959 = ((~g10402));
assign g11049 = ((~II16808));
assign g4069 = (g1762&g2802);
assign g2938 = ((~II6110))|((~II6111));
assign g7675 = ((~II12300));
assign g9335 = (g8975&g5708);
assign g3281 = (g766&g2525);
assign g4000 = (g1744&g2778);
assign g5194 = (g1610&g4717);
assign g8687 = (g8558&g8036);
assign g6819 = (g243&g6596);
assign g6563 = ((~g5783));
assign II6761 = ((~g2943))|((~II6760));
assign g4995 = (g1474&g4640);
assign g3062 = ((~g2369))|((~g591))|((~g611));
assign g8307 = ((~II13294))|((~II13295));
assign g9389 = (g1330&g9151);
assign g6360 = (g302&g5899);
assign II5751 = ((~g2296));
assign g10357 = (g10278&g2462);
assign II16514 = ((~g10717));
assign g5024 = (g1284&g4513);
assign g8968 = (g8089&g6778&g8849);
assign II7691 = ((~g3363));
assign g10179 = ((~g10041));
assign II14866 = (g9590)|(g9609)|(g9619);
assign g9900 = (g9845&g8327);
assign g7892 = (g7616&g3815);
assign II7684 = ((~g1023))|((~II7683));
assign g3774 = ((~II6999));
assign II10141 = ((~g5683));
assign g9907 = (g9888&g9686);
assign g7089 = ((~II11322));
assign II4894 = ((~g258));
assign II7683 = ((~g1023))|((~g3460));
assign II14525 = ((~g9109));
assign g4355 = ((~II7642));
assign g7026 = ((~II11173));
assign g8447 = ((~II13639));
assign g4610 = (g3804&g2212);
assign g4940 = (g3500&g4440);
assign II7375 = ((~g4062));
assign g4396 = ((~II7735));
assign g6365 = ((~II10274));
assign g10195 = ((~II15559));
assign II12128 = ((~g170))|((~II12126));
assign g8191 = ((~II13114));
assign g7982 = ((~II12790));
assign g10042 = ((~II15253));
assign g3412 = (g219&g3228);
assign II6501 = ((~g2578));
assign g8995 = (g6454&g8929);
assign II13300 = ((~g1936))|((~g8162));
assign g3436 = ((~g3144));
assign II6331 = (g2060&g2070&g2074&g2077);
assign II7381 = ((~g4078));
assign II6827 = ((~g770))|((~II6825));
assign g6542 = (g5789)|(g5010);
assign g7763 = ((~II12454));
assign g9569 = (g9052)|(g9030);
assign g10535 = ((~II16172));
assign II17347 = ((~g11373));
assign g4556 = (g3536)|(g2916);
assign II10849 = ((~g6734));
assign g5729 = ((~II9279));
assign II5513 = ((~g255));
assign II15400 = ((~g10069));
assign g2368 = ((~II5445));
assign g6561 = ((~g5773));
assign g4311 = ((~g4130));
assign g6293 = ((~II10138));
assign g5788 = (g1540&g5231);
assign g11249 = (g6162)|(g11143);
assign g11061 = ((~g10974));
assign g11238 = (g5474&g11110);
assign g6577 = ((~II10520))|((~II10521));
assign g7911 = ((~g7664));
assign g6201 = ((~II9938));
assign II6106 = ((~g2116));
assign g5748 = ((~II9320));
assign g11305 = (g11215)|(g11093);
assign g5805 = ((~II9409));
assign g5216 = ((~g4445));
assign g11467 = ((~II17438));
assign g7352 = ((~II11704));
assign g11092 = (g837&g10950);
assign g6629 = ((~II10584));
assign g5025 = (g1482&g4640);
assign II16607 = ((~g10787));
assign g7314 = ((~II11590));
assign g10913 = ((~II16691));
assign g2098 = ((~II4938));
assign II17202 = ((~g11322));
assign g10571 = ((~II16236));
assign g9785 = (g9010)|(g8995)|(g9388)|(g9363);
assign g2455 = ((~g826));
assign g4342 = (g1149&g3719);
assign II17758 = ((~g11647));
assign g5445 = (g4631&g3875&g2733);
assign g4432 = (g3723&g1975);
assign g3761 = ((~II6962));
assign g8361 = ((~II13463));
assign g7367 = (g7224)|(g6744);
assign II7999 = ((~g4114));
assign g5680 = (g153&g5361);
assign g4835 = ((~II8192));
assign g7030 = ((~II11183));
assign g4197 = ((~II7408));
assign g10666 = (g10575&g9424);
assign II13661 = ((~g8322))|((~II13659));
assign II17121 = ((~g11231));
assign g6419 = ((~II10331));
assign g7696 = ((~g7148));
assign g8319 = ((~II13341));
assign g10561 = (g10549&g4583);
assign g11325 = (g11295)|(g11165);
assign g8892 = ((~II14242));
assign g6261 = ((~II10042));
assign II5722 = ((~g2075));
assign g8728 = (g8610&g7915);
assign g4009 = (g1747&g2789);
assign II14786 = ((~g9266));
assign g2859 = ((~II5995));
assign g4236 = (g1098&g3638);
assign g9715 = (g1531&g9490);
assign II11804 = ((~g7190));
assign g8532 = ((~II13741));
assign g10174 = ((~II15514));
assign g8403 = (g6101&g8239);
assign II6208 = ((~g2534))|((~II6207));
assign II16571 = ((~g10819));
assign g3119 = ((~II6347));
assign g6872 = (g1896&g6389);
assign g2298 = ((~II5336));
assign g5498 = ((~II8919));
assign g5874 = ((~II9491));
assign g10550 = (g4942)|(g10450);
assign II5185 = ((~g1415))|((~II5184));
assign g4401 = (g2971&g3772);
assign II9973 = ((~g5502));
assign g9879 = ((~g9747)&(~g9536)&(~g9566)&(~II15048));
assign g7214 = ((~II11450));
assign g8119 = (g6239&g7890);
assign II5957 = ((~g2178));
assign g8170 = (g5270&g7853);
assign II12556 = ((~g7678));
assign II9673 = ((~g5182));
assign II14862 = (g9587)|(g9600)|(g9611);
assign II8529 = ((~g481))|((~II8527));
assign g7604 = ((~II12162));
assign g7073 = ((~II11296));
assign g4454 = ((~g3914));
assign g11424 = ((~II17327));
assign g3474 = ((~II6679));
assign g8780 = ((~II14077));
assign g10349 = ((~II15811));
assign g10417 = (g10301)|(g9527);
assign II12144 = ((~g7089))|((~II12143));
assign g7192 = ((~g6742));
assign II16295 = ((~g10552));
assign g6853 = ((~II10917));
assign g8749 = (g7604&g8660);
assign g9594 = (g1&g9292);
assign g7064 = ((~II11269));
assign g4212 = ((~II7453));
assign g4811 = ((~g3661));
assign g10176 = ((~II15520));
assign g8779 = (g5530)|(g8663);
assign II12907 = ((~g7959));
assign g7457 = (g6873)|(g6404);
assign g5983 = (g5084)|(g4392);
assign II15798 = ((~g10281));
assign g9849 = (g293&g9768);
assign g8314 = ((~II13326));
assign g3067 = ((~II6273));
assign II7606 = ((~g4166));
assign II9769 = ((~g5287));
assign g4421 = (g4112&g2980);
assign g6879 = (g1914&g6407);
assign g7895 = (g7503&g7036);
assign II15205 = (g9838)|(g9963)|(g9850)|(g9878);
assign g10681 = (g10567&g3586);
assign g6837 = ((~II10891));
assign g3716 = ((~II6876));
assign g5743 = ((~II9311));
assign II7651 = ((~g3332));
assign II15418 = ((~g10083));
assign g8075 = (g727&g7826);
assign g11437 = ((~II17362));
assign g7626 = (g7060)|(g5267);
assign g3404 = ((~g3121));
assign g6923 = (g6353)|(g5695);
assign II17704 = ((~g11618));
assign II6013 = ((~g2200));
assign g10784 = (g10727&g5169);
assign g6942 = ((~II11076));
assign g5694 = (g162&g5361);
assign II10974 = ((~g6563));
assign II11599 = ((~g6832));
assign g6994 = (g6758&g3829);
assign g7450 = ((~g7148));
assign g2018 = ((~g1336));
assign g9767 = ((~II14914));
assign g8385 = (g6084&g8218);
assign g6587 = ((~g5827));
assign g7938 = ((~g7403));
assign II16641 = ((~g10864));
assign g7523 = ((~II11908))|((~II11909));
assign II15250 = ((~g9980));
assign II6941 = ((~g2858));
assign g6549 = (g5515&g6175);
assign II13515 = ((~g8248))|((~II13513));
assign II10807 = ((~g6396));
assign g6523 = (g5745)|(g4995);
assign II12199 = ((~g7278));
assign g4068 = (g2719&g2276);
assign g4419 = ((~II7763));
assign g4526 = ((~II7931));
assign g4144 = ((~g2160))|((~g3044));
assign g8757 = ((~g8599))|((~g4401));
assign g4619 = ((~g3077)&(~g3491)&(~g3485)&(~g2655));
assign g11595 = (g1336&g11575);
assign g8520 = ((~II13729));
assign II8787 = ((~g4639))|((~II8786));
assign II15956 = ((~g10402));
assign II8358 = ((~g4794));
assign g4481 = (g1713&g3906);
assign g3333 = ((~g2779));
assign g4114 = (g1351&g3301);
assign g4756 = ((~g3440));
assign g6556 = ((~g5747));
assign g11514 = (g11491&g5151);
assign II13200 = ((~g8251));
assign g3010 = ((~g2382))|((~g2399));
assign II14005 = ((~g8631));
assign g5758 = ((~II9338));
assign II8652 = ((~g778))|((~II8650));
assign g5478 = (g1905&g4242);
assign II5174 = ((~g52));
assign g4839 = (g225&g3946);
assign g4208 = ((~II7441));
assign g3438 = (g2939)|(g2944);
assign II10685 = ((~g6054));
assign g11034 = ((~II16763));
assign g6951 = ((~II11097));
assign II5690 = (g1436&g1440&g1444&g1448);
assign II14573 = ((~g9029));
assign g7936 = ((~g7712));
assign g10625 = (g10546&g4552);
assign g2833 = ((~II5949));
assign II17719 = ((~g11623));
assign II13027 = ((~g8051));
assign g6396 = ((~II10296));
assign g7991 = ((~II12809));
assign II17770 = ((~g11649));
assign g11507 = ((~II17540));
assign g9764 = ((~g9432));
assign II13194 = ((~g8140));
assign g2547 = ((~g23));
assign II15033 = (g7853)|(g9804)|(g9624)|(g9785);
assign g6208 = ((~II9953));
assign g8787 = ((~II14094));
assign g7677 = ((~g7148));
assign g5814 = (g5591)|(g4827);
assign g10342 = ((~II15792));
assign II16387 = ((~g10629));
assign II16656 = ((~g10791));
assign g11009 = (g5179&g10827);
assign II7086 = ((~g3142));
assign II17505 = ((~g7603))|((~II17503));
assign g7045 = ((~g6435));
assign II9221 = ((~g5236));
assign II11275 = ((~g6502));
assign g3399 = (g2918)|(g2940);
assign II5014 = ((~g1007))|((~II5013));
assign g4178 = ((~II7351));
assign g3768 = ((~II6979));
assign g7023 = ((~II11166));
assign II14873 = ((~g9525));
assign II10322 = ((~g6193));
assign g11357 = ((~II17182));
assign g3382 = ((~II6580));
assign g5541 = (g4331&g3582);
assign g5198 = ((~II8614));
assign II10639 = ((~g5830));
assign g3912 = (g207&g3164);
assign II6360 = ((~g2261));
assign II9458 = ((~g5091));
assign g10374 = ((~g10347)&(~g3463));
assign g8680 = ((~II13965));
assign g10366 = ((~g10285))|((~g5392));
assign g9384 = (g968&g9223);
assign g2356 = ((~II5438));
assign g5269 = ((~II8716))|((~II8717));
assign g8766 = (g8612&g5151);
assign II16269 = ((~g10558));
assign g5629 = ((~II9065));
assign g9028 = ((~II14421));
assign g6055 = ((~II9688));
assign II16518 = ((~g10718));
assign g4266 = ((~g3688));
assign g2078 = ((~g135));
assign g8986 = ((~II14379));
assign g2915 = ((~II6094));
assign g9560 = (g9052)|(g9030);
assign g9750 = ((~g9454)&(~g9274)&(~g9292));
assign II7423 = ((~g3331));
assign II8388 = ((~g4239));
assign g4542 = (g366&g3586);
assign g7539 = ((~II11953));
assign g10320 = ((~II15756));
assign g9317 = (g6109&g8875);
assign g8558 = ((~II13766))|((~II13767));
assign g2112 = ((~g639));
assign II16142 = (g10511&g10509&g10507);
assign g4603 = ((~g3829));
assign g6093 = (g5264)|(g4534);
assign g6185 = (g5470)|(g4715);
assign II15225 = (g9842)|(g9967)|(g9859)|(g9881);
assign g7219 = (g6661)|(g6076);
assign g1983 = ((~g750));
assign II10355 = ((~g6003));
assign g4207 = ((~II7438));
assign II11814 = ((~g7196));
assign g8051 = (g7572&g5128);
assign g9951 = (g9902)|(g9899)|(g9803);
assign II13469 = ((~g8147));
assign g11401 = ((~II17246));
assign g7925 = ((~g7476));
assign II14370 = ((~g8954));
assign g5047 = ((~g4354));
assign II14964 = ((~g9762));
assign g10286 = ((~g10271)&(~g3463));
assign II6792 = ((~g2959))|((~g143));
assign g3003 = ((~g599))|((~g2399));
assign g10254 = ((~g10196));
assign g5916 = ((~II9550));
assign g10471 = ((~g10378));
assign g11469 = ((~II17444));
assign g8186 = ((~II13109));
assign g2796 = ((~g2276));
assign g5536 = (g4867&g4298);
assign II11029 = ((~g6485));
assign g7321 = ((~II11611));
assign g2389 = ((~II5469))|((~II5470));
assign II7889 = ((~g3373));
assign g5396 = (g4481)|(g3684);
assign g7996 = ((~g7011))|((~g7574))|((~g7562))|((~g6974));
assign g4803 = ((~g3664))|((~g2356));
assign II15608 = ((~g10149))|((~II15607));
assign g3094 = ((~II6302));
assign g6239 = ((~II9988));
assign g4333 = ((~g4144));
assign II17586 = ((~g11515))|((~II17584));
assign II10240 = ((~g5937));
assign g2534 = (g798&g794);
assign g3400 = (g115&g3164);
assign II6965 = ((~g2880));
assign II5101 = ((~g1960));
assign g11540 = ((~g11519));
assign g11620 = ((~II17678));
assign g8324 = ((~II13354));
assign g9515 = (g9173)|(g9151);
assign g9872 = (g9617)|(g9594)|(g9750);
assign II17519 = ((~g11484));
assign II11647 = ((~g6925));
assign g4294 = ((~g3664));
assign g8045 = (g7547&g5128);
assign g7784 = ((~II12517));
assign g3077 = ((~g2213));
assign g9410 = ((~g9010)&(~g9240)&(~g9223)&(~II14607));
assign II13442 = ((~g8182));
assign g8750 = ((~II14045));
assign g9361 = ((~g9010)&(~g9240)&(~g9223)&(~II14582));
assign II9380 = ((~g5013));
assign g3772 = (g2542&g3089);
assign g2419 = ((~II5501))|((~II5502));
assign II17724 = ((~g11625));
assign II15906 = ((~g6899))|((~g10302));
assign II8543 = ((~g4218))|((~g486));
assign II6282 = ((~g2231));
assign g10499 = ((~II16124));
assign II10099 = ((~g5800));
assign g11168 = (g534&g11112);
assign g8340 = ((~II13400));
assign g8004 = ((~II12838));
assign g11014 = ((~II16735));
assign II12871 = ((~g7638));
assign g2450 = ((~g1351));
assign g2561 = (g742&g741);
assign II5166 = ((~g1499))|((~II5164));
assign g3329 = ((~II6504));
assign g7680 = ((~g7148));
assign II13475 = ((~g8173));
assign g11558 = (g2713&g11519);
assign g8479 = ((~g8319));
assign II14914 = ((~g9533));
assign g4566 = ((~g3753));
assign II16720 = ((~g10854));
assign g11440 = ((~II17371));
assign g2847 = ((~II5973));
assign II12086 = ((~g6980))|((~II12085));
assign II8797 = ((~g1145))|((~II8795));
assign II15688 = ((~g10207));
assign g6857 = ((~II10927));
assign g7725 = ((~II12360));
assign g9935 = (g9914&g9624);
assign g8033 = ((~II12875));
assign g11430 = (g11387)|(g4006);
assign g4880 = ((~g3638));
assign II10302 = ((~g6179));
assign g6327 = (g1255&g5949);
assign II9062 = ((~g4759));
assign g5548 = ((~g1840))|((~g4401));
assign g5601 = (g1035&g4375);
assign g10686 = (g10612&g3863);
assign g2719 = ((~g2043));
assign g9701 = (g1574&g9474);
assign g10523 = ((~g10456));
assign II14827 = (g9603)|(g9614)|(g9584);
assign g6434 = ((~II10352));
assign g4002 = ((~g3121));
assign g5527 = ((~g3978))|((~g4749));
assign g10698 = ((~II16373));
assign II8606 = ((~g506))|((~II8604));
assign g9644 = (g1182&g9125);
assign g4012 = ((~II7154));
assign g8876 = (g8105&g6764&g8858);
assign g7202 = (g6349&g4329);
assign g9583 = (g886&g8995);
assign II12469 = ((~g7531));
assign II6028 = ((~g2208));
assign II17216 = ((~g11291));
assign II13868 = ((~g8523))|((~II13867));
assign g8064 = ((~II12910));
assign g2082 = ((~g1371));
assign g7379 = ((~g6863));
assign g10395 = ((~g10320));
assign g11649 = ((~II17749));
assign g5948 = ((~II9588));
assign g7817 = ((~II12616));
assign g2961 = ((~II6177))|((~II6178));
assign II7408 = ((~g4125));
assign II16760 = ((~g10888));
assign II5529 = ((~g1265))|((~II5528));
assign g10578 = ((~g10527));
assign g8168 = (g5262&g7853);
assign g11052 = ((~II16817));
assign II9836 = ((~g5405));
assign II10941 = ((~g6555));
assign g4387 = ((~II7716));
assign g10309 = ((~II15733));
assign g6301 = ((~II10162));
assign II16114 = ((~g10387));
assign g5996 = (g5473)|(g3908);
assign II12137 = ((~g7110))|((~II12136));
assign g5191 = ((~g4640));
assign g6197 = ((~II9930));
assign II12502 = ((~g7726));
assign II14194 = ((~g8798));
assign g11389 = ((~II17216));
assign g9597 = (g1170&g9125);
assign g5203 = ((~g4640));
assign g11273 = (g5638&g11195);
assign g4900 = ((~II8265));
assign II16897 = ((~g10947));
assign g2980 = ((~g1983));
assign II5538 = ((~g1270))|((~g1023));
assign g4259 = ((~g3292)&(~g3793)&(~g3784)&(~g3776));
assign g7328 = ((~II11632));
assign g11441 = ((~II17374));
assign g8302 = ((~II13273))|((~II13274));
assign g2248 = ((~g99));
assign g4076 = ((~g1707)&(~g2864));
assign g10726 = (g10316)|(g10673);
assign II6985 = ((~g2890));
assign II6201 = ((~g766))|((~II6199));
assign g5177 = ((~g4596));
assign g11419 = ((~II17312));
assign g7055 = (g5900&g6579);
assign II15395 = ((~g10058));
assign g8246 = (g7846&g7442);
assign g3506 = (g986&g2760);
assign g5040 = ((~II8421));
assign g8716 = ((~g8576));
assign g10881 = ((~II16613));
assign II11243 = ((~g790))|((~II11241));
assign g2515 = ((~II5605))|((~II5606));
assign g6226 = ((~II9973));
assign II13227 = ((~g8264));
assign g11310 = (g11220)|(g11100);
assign g8355 = ((~II13445));
assign g9808 = ((~g9392)&(~g9367));
assign g5676 = ((~II9185));
assign II5378 = ((~g1857));
assign g4382 = ((~g3638));
assign II8738 = ((~g4607))|((~g1121));
assign g2850 = ((~II5976));
assign g11486 = (g6654)|(g11463);
assign g9926 = (g9868)|(g9715);
assign II10374 = ((~g5852));
assign g10450 = (g10364&g3359);
assign g4225 = ((~II7478));
assign g4565 = (g534&g4010);
assign g4188 = ((~II7381));
assign II12933 = ((~g7899));
assign g2606 = ((~II5719));
assign g7052 = ((~II11235));
assign g7568 = ((~II12026));
assign II14697 = ((~g9260));
assign g8245 = (g7850&g4339);
assign g3661 = (g382&g3257);
assign g5421 = (g4631&g2733&g3819);
assign g6420 = ((~II10334));
assign g7093 = ((~II11326));
assign g4222 = ((~g3638));
assign II13639 = ((~g8321));
assign II17675 = ((~g11606));
assign g5687 = (g139&g5361);
assign g11609 = (g11588)|(g11559);
assign II12641 = ((~g7709));
assign g10231 = ((~II15616))|((~II15617));
assign g2126 = ((~g12));
assign g3829 = (g2028&g2728);
assign g4607 = ((~g3077)&(~g2669)&(~g3485)&(~g3479));
assign II11829 = ((~g7213));
assign II7143 = ((~g2614));
assign II9282 = ((~g5633));
assign II17053 = ((~g11249))|((~II17051));
assign g11185 = ((~II16956));
assign g10158 = ((~II15470));
assign g2116 = ((~II5020));
assign g9953 = (g9945)|(g9939)|(g9669);
assign II15756 = ((~g10266));
assign II16879 = ((~g10936));
assign g8068 = (g664&g7826);
assign g6214 = ((~g5446));
assign g7821 = (g1905&g7479);
assign g10638 = (g10608&g3829);
assign II10623 = ((~g6002));
assign g6444 = ((~g6158));
assign II7843 = ((~g3440));
assign II17610 = ((~g11549));
assign g7069 = ((~II11286));
assign g9261 = ((~g8892));
assign g6355 = ((~g6032)&(~g6023));
assign g9619 = (g2772&g9010);
assign g5004 = (g1296&g4499);
assign g5797 = ((~II9399));
assign g10474 = ((~II16024))|((~II16025));
assign g2091 = (g976&g971);
assign g10731 = (g5118&g1850&g10665);
assign II7191 = ((~g2646));
assign II12076 = ((~g174))|((~II12074));
assign II11188 = ((~g6513));
assign g5085 = ((~g4377));
assign g10448 = (g10421&g3335);
assign g5515 = ((~g4429));
assign g4061 = ((~II7182));
assign II7735 = ((~g3759));
assign II10560 = ((~g5887));
assign g2343 = ((~g1927));
assign g8470 = (g8308&g7427);
assign g4096 = ((~II7236));
assign g5617 = (g1050&g4391);
assign II13295 = ((~g8161))|((~II13293));
assign g9424 = ((~g9076));
assign II7112 = ((~g3186));
assign g8823 = (g8778)|(g8693);
assign g8970 = ((~g5548))|((~g8839));
assign II15244 = ((~g10031));
assign g8412 = ((~II13545))|((~II13546));
assign g8349 = ((~II13427));
assign g11208 = ((~g11077));
assign II7321 = ((~g3047))|((~g1231));
assign II10573 = ((~g5980));
assign II13460 = ((~g8155));
assign g3684 = (g1710&g3015);
assign II5815 = ((~g1994));
assign II13323 = ((~g8203));
assign g7905 = ((~g7450));
assign II11263 = ((~g826))|((~II11261));
assign g10871 = ((~II16583));
assign g4585 = (g521&g4060);
assign g10467 = ((~II15993))|((~II15994));
assign g4180 = ((~II7357));
assign g3253 = ((~II6417));
assign g10878 = ((~II16604));
assign II13090 = ((~g8006))|((~II13089));
assign g3290 = ((~II6461));
assign g2438 = ((~g243));
assign II12388 = ((~g7219));
assign g4502 = (g2031&g3938);
assign g9708 = (g9653)|(g9389)|(g9646);
assign II8406 = ((~g4274));
assign II6196 = ((~g2462));
assign g6044 = ((~II9665));
assign g5846 = (g4932)|(g4236);
assign II6468 = ((~g23))|((~II6467));
assign g9603 = (g1173&g9125);
assign II5809 = ((~g2356));
assign II17084 = ((~g11249));
assign g6616 = (g6105&g3246);
assign g2906 = ((~II6071));
assign g11642 = ((~II17730));
assign g2754 = ((~II5830));
assign II10831 = ((~g6710));
assign g3782 = ((~II7006));
assign II17558 = ((~g11504));
assign II10508 = ((~g6221))|((~II10507));
assign g2613 = ((~II5740));
assign II11071 = ((~g6656));
assign II12759 = ((~g7702));
assign II5684 = ((~g572));
assign g5937 = ((~II9567));
assign g2601 = ((~II5704));
assign g2243 = ((~II5248));
assign g4954 = ((~g4509));
assign II9953 = ((~g5484));
assign g10851 = ((~II16553));
assign II6226 = ((~g1346))|((~II6224));
assign g9909 = (g9891&g9804);
assign g5492 = (g1654&g4263);
assign II9174 = ((~g4903));
assign g11191 = ((~g11112));
assign g6812 = ((~II10846));
assign g2608 = ((~II5725));
assign II5254 = ((~g1700));
assign g2626 = ((~g2000));
assign g7635 = ((~II12245));
assign g9831 = (g9727&g9785);
assign g3106 = ((~II6323))|((~II6324));
assign II12862 = ((~g7638));
assign g6102 = (g1038&g5320);
assign g9718 = (g1540&g9490);
assign g11471 = ((~II17450));
assign g4103 = (g2683&g2997);
assign g2179 = ((~g89));
assign g9728 = (g9412)|(g9422)|(g9426);
assign II16413 = ((~g10663));
assign g6828 = (g1377&g6596);
assign g10684 = (g10604&g3863);
assign g4723 = (g3626&g2779);
assign II9779 = ((~g5391));
assign g11231 = (g11156)|(g11013);
assign g10518 = (g10513&g10440&II16145);
assign g2158 = ((~II5077));
assign II5383 = ((~g886));
assign g11474 = ((~II17460))|((~II17461));
assign g2104 = ((~II4965))|((~II4966));
assign g11546 = ((~g11519));
assign II11767 = ((~g7201));
assign II12087 = ((~g1470))|((~II12085));
assign g6817 = ((~II10861));
assign g8144 = ((~II13027));
assign g8516 = ((~II13717));
assign g4451 = ((~g3638));
assign g5499 = (g1627&g4270);
assign g5009 = (g1486&g4640);
assign g6535 = (g345&g6063);
assign g7650 = ((~II12261));
assign g11016 = ((~II16739));
assign II10873 = ((~g6331));
assign g9961 = ((~II15162));
assign g8972 = (g8085&g6764&g8858);
assign g2184 = ((~g1806));
assign g5319 = ((~II8804))|((~II8805));
assign g9940 = (g9920&g9367);
assign g11111 = ((~g10974));
assign II12487 = ((~g7723));
assign g7943 = (g2840&g7467);
assign II10251 = ((~g6126));
assign II11904 = ((~g6902));
assign g6111 = ((~II9786));
assign g9447 = (g1762&g9030);
assign II12986 = ((~g8042));
assign II6748 = ((~g1453))|((~II6746));
assign g8646 = (g8224)|(g8547);
assign g2800 = (g2399&g2369&g591);
assign g8507 = ((~g3738))|((~g8366));
assign g4991 = (g1508&g4640);
assign II9243 = ((~g5245));
assign II9829 = ((~g5013));
assign g4291 = ((~g4013));
assign g9354 = ((~II14567));
assign g10318 = ((~II15752));
assign g10929 = ((~g10827));
assign II7444 = ((~g3683));
assign g3743 = ((~II6932));
assign g6135 = ((~II9842));
assign g6543 = ((~g5888));
assign g4063 = (g2713&g2276);
assign g7562 = ((~g6984));
assign II15771 = ((~g10250));
assign II17633 = ((~g11578));
assign g7243 = ((~II11483));
assign g8118 = (g1900&g7941);
assign g7571 = ((~II12035));
assign g8703 = (g7601&g8585);
assign g4156 = ((~II7295));
assign g11643 = ((~II17733));
assign g4961 = ((~II8333));
assign II15548 = ((~g10083));
assign g9622 = (g1200&g9111);
assign g7556 = ((~II11992));
assign g11144 = (g305&g10926);
assign g2199 = ((~g48));
assign g7804 = ((~II12577));
assign II11159 = ((~g6478));
assign g11215 = (g953&g11160);
assign g4479 = ((~II7858));
assign g8651 = (g8520&g4013);
assign g7606 = ((~II12168));
assign g3379 = ((~g3121));
assign g6427 = ((~II10343));
assign II5308 = ((~g97));
assign II15458 = ((~g10069));
assign II8804 = ((~g4677))|((~II8803));
assign g5914 = (g5029)|(g4343);
assign g6500 = (g5725)|(g4986);
assign g5250 = (g1270&g4748);
assign g6697 = ((~g5949));
assign gbuf4 = (g874);
assign II9717 = ((~g5426));
assign II10584 = ((~g5864));
assign g9902 = (g9894&g9392);
assign g10482 = ((~II16080))|((~II16081));
assign g10742 = (g10655&g3586);
assign g1993 = ((~g786));
assign g5777 = ((~II9365));
assign g7508 = ((~g6950));
assign II9655 = ((~g5173));
assign g3220 = ((~II6398));
assign II17485 = ((~g11384))|((~g11474));
assign g8981 = ((~II14364));
assign II14340 = ((~g8820));
assign g6896 = ((~II10996));
assign II9402 = ((~g5107));
assign g9474 = ((~g9331));
assign g10485 = (g9317)|(g10376);
assign g5608 = (g814&g4831);
assign II6546 = ((~g2987));
assign g8261 = (g7876)|(g3383);
assign II15804 = ((~g10283));
assign g8287 = (g8117)|(g7824);
assign g6271 = ((~II10072));
assign g6350 = (g5837&g4435);
assign g2844 = ((~II5966));
assign II5104 = ((~g431))|((~g435));
assign II12913 = ((~g7845));
assign II16947 = ((~g11080));
assign g8642 = (g5236)|(g5205)|(g8465);
assign g7757 = ((~II12436));
assign g8975 = (g8089&g6764&g8858);
assign g9605 = ((~g9125)&(~g9111)&(~g9173)&(~g9151));
assign g10753 = (g10649&g4013);
assign g8469 = (g8305&g7422);
assign II7771 = ((~g3418));
assign g8462 = (g8300&g7406);
assign II12251 = ((~g7076));
assign II6136 = ((~g2496))|((~g378));
assign g10311 = ((~g10242));
assign g9363 = (g9205)|(g9192);
assign g8053 = (g7583&g5919);
assign g11343 = ((~II17152));
assign II14270 = ((~g8840))|((~g1822));
assign g4057 = ((~II7176));
assign g10133 = ((~g10064));
assign II11534 = ((~g6917));
assign g4898 = ((~II8259));
assign g7505 = ((~g7148));
assign g9869 = (g1558&g9814);
assign II12177 = ((~g7259));
assign II8780 = ((~g1137))|((~II8778));
assign g8940 = (g8793)|(g8703);
assign g11031 = (g411&g10974);
assign g9695 = (g1567&g9474);
assign II11701 = ((~g7065));
assign II7563 = ((~g3533))|((~II7562));
assign g4460 = ((~g3820));
assign II13648 = ((~g8376));
assign II8561 = ((~g4227))|((~g491));
assign II17283 = ((~g11357))|((~II17281));
assign g7589 = ((~II12099));
assign g3696 = (g1713&g3015);
assign g10669 = (g10577&g9429);
assign g6268 = ((~II10063));
assign g5936 = ((~II9564));
assign g10765 = (g5492)|(g10680);
assign g6663 = (g6064&g2237);
assign II13373 = ((~g8226));
assign II14349 = ((~g8958));
assign g4160 = ((~II7303));
assign g4998 = (g1304&g4485);
assign g4932 = (g1065&g4442);
assign II13412 = ((~g8142));
assign II5707 = ((~g2418));
assign II11312 = ((~g6488));
assign g7289 = ((~II11543));
assign g8239 = ((~g7826));
assign g6125 = ((~II9822));
assign g6748 = ((~II10753));
assign g5006 = (g1462&g4640);
assign g8010 = (g7738&g7413);
assign g2701 = ((~g2040));
assign g8164 = ((~g7872));
assign II15451 = ((~g10058))|((~g10051));
assign g2839 = ((~II5957));
assign g9432 = ((~g9313));
assign II15323 = ((~g10019));
assign g5106 = ((~II8490));
assign II13747 = ((~g8299));
assign g2015 = ((~g1107));
assign II6870 = ((~g2852));
assign g4218 = ((~g3292)&(~g2593)&(~g3784)&(~g3776));
assign g9610 = (g925&g9192);
assign g8555 = (g8409&g8025);
assign II17374 = ((~g11411));
assign g4374 = ((~II7684))|((~II7685));
assign g9573 = (g9052)|(g9030);
assign II14185 = ((~g8790));
assign g8172 = (g5275&g7853);
assign g8138 = ((~II13013));
assign g4675 = ((~g4073))|((~g3247));
assign g11634 = ((~II17716));
assign II9093 = ((~g5397));
assign g11617 = ((~II17669));
assign g7290 = (g7046)|(g6316);
assign II9798 = ((~g5415));
assign g7536 = (g7148&g2877);
assign g11154 = (g330&g10932);
assign g2329 = ((~II5383));
assign g6738 = (g2531&g6137);
assign g8884 = ((~II14224));
assign g4778 = (g421&g3426);
assign II11037 = ((~g6629));
assign II15377 = ((~g10104));
assign II16867 = ((~g10913));
assign II16592 = ((~g10781));
assign II9156 = ((~g5032));
assign II10243 = ((~g5918));
assign g6334 = (g1389&g5904);
assign g4865 = (g1080&g3638);
assign g6755 = (g6106)|(g5479);
assign II9783 = ((~g5395));
assign g8383 = (g8163)|(g5051);
assign g11585 = (g1321&g11543);
assign g3683 = ((~II6844));
assign g9739 = ((~II14884));
assign g8437 = ((~II13609));
assign g10559 = (g4141)|(g10512);
assign g6744 = (g4828&g6151);
assign g7657 = ((~II12268));
assign g2550 = ((~g1834));
assign II6639 = ((~g2632));
assign g4716 = ((~g3546));
assign g8025 = ((~II12867));
assign g6363 = (g284&g5901);
assign g5660 = ((~II9141));
assign g11339 = ((~II17142));
assign g8500 = ((~II13695));
assign g8105 = ((~g7992));
assign g10496 = (g10429&g3977);
assign II8772 = ((~g1133))|((~II8770));
assign g9240 = (g6454&g8962);
assign II8795 = ((~g4672))|((~g1145));
assign g9646 = ((~g9125)&(~g9151));
assign II17470 = ((~g11452));
assign g7135 = (g869&g6355);
assign II8664 = ((~g476))|((~II8662));
assign g6035 = (g5518)|(g3974);
assign II14543 = ((~g9311));
assign II5399 = ((~g895));
assign g7595 = ((~II12123));
assign g10114 = ((~II15350));
assign g7298 = (g7136)|(g6324);
assign II7648 = ((~g3727));
assign II5084 = (g1462&g1470&g1474&g1478);
assign g5186 = ((~g2047)&(~g4401));
assign g9680 = (g9454)|(g9292)|(g9274);
assign II9032 = ((~g4732));
assign g10490 = ((~II16105));
assign g4884 = (g3813&g2971);
assign g4126 = (g2701&g3040);
assign g7729 = ((~II12372));
assign II8996 = ((~g4757));
assign g8807 = ((~II14140));
assign g7131 = (g6044&g6700);
assign g7796 = ((~II12553));
assign g5981 = (g5074)|(g4383);
assign g1988 = ((~g766));
assign g2726 = ((~g2021));
assign g4966 = ((~II8340));
assign g10782 = (g10725&g5146);
assign g11574 = ((~g11561));
assign II5451 = ((~g991))|((~II5449));
assign g2252 = ((~II5271));
assign g10334 = (g10265&g3307);
assign g5253 = ((~g4346));
assign g5943 = ((~II9581));
assign II12061 = ((~g6961))|((~II12060));
assign g10923 = (g10778)|(g10715);
assign g6310 = ((~II10189));
assign II8839 = ((~g4484));
assign g9913 = (g9849)|(g9691);
assign g4414 = ((~II7752));
assign g9964 = (g9954&g9536);
assign II15586 = ((~g10159));
assign g7237 = ((~II11477));
assign g8736 = (g7439&g8635);
assign g6507 = (g5732)|(g4990);
assign II4917 = ((~g584));
assign g10893 = ((~II16641));
assign II6664 = ((~g2792))|((~g2776));
assign II14596 = (g8995)|(g9205)|(g9192);
assign g10793 = (g6194)|(g10763);
assign II5731 = ((~g2089));
assign g6156 = ((~g5426));
assign g6141 = ((~II9854));
assign II5501 = ((~g1255))|((~II5500));
assign g7230 = (g6064&g6444);
assign g6236 = ((~II9981));
assign II13720 = ((~g8358));
assign II9409 = ((~g5013));
assign g11492 = (g11480&g4807);
assign g7615 = ((~II12193));
assign g8663 = (g8538&g4013);
assign g2882 = ((~II6034));
assign g7592 = ((~II12107))|((~II12108));
assign II6166 = ((~g2236))|((~g153));
assign g3704 = ((~II6861));
assign II14681 = ((~g9110));
assign g7662 = ((~II12279));
assign II10461 = ((~g5849));
assign II16079 = ((~g849))|((~g10374));
assign g4047 = (g2695&g2276);
assign II14352 = ((~g8946));
assign g9125 = (g8966&g6674);
assign g2372 = ((~II5450))|((~II5451));
assign g4733 = ((~II8089));
assign g6219 = ((~g5426));
assign II13114 = ((~g7930));
assign g7669 = ((~II12286));
assign g11456 = (g3765&g3517&g11422);
assign II6513 = ((~g2812));
assign II6802 = ((~g2751));
assign II10655 = ((~g6036));
assign g2202 = ((~g148));
assign II11964 = ((~g6910));
assign II15335 = ((~g10007));
assign g10504 = (g10389&g2135);
assign g4821 = ((~II8179))|((~II8180));
assign g5863 = (g5272&g2173);
assign g6417 = ((~g6136));
assign g11088 = ((~II16871));
assign g7971 = (g5110)|(g7549);
assign g3326 = ((~II6495));
assign g2335 = ((~II5391));
assign II10054 = ((~g5728));
assign g7148 = ((~II11397));
assign g8630 = ((~II13908))|((~II13909));
assign II11740 = ((~g7030));
assign II5737 = ((~g2100));
assign g6144 = ((~II9857));
assign g4682 = (g3563)|(g3348)|(g1570);
assign g7786 = ((~II12523));
assign II8670 = ((~g4831))|((~II8669));
assign II13794 = ((~g8472));
assign g2042 = ((~g1796));
assign g8036 = ((~II12878));
assign II12021 = ((~g166))|((~II12019));
assign g10164 = ((~II15488));
assign g10383 = ((~g10318)&(~g2998));
assign II17164 = ((~g11320));
assign II15045 = (g7853)|(g9676)|(g9624)|(g9785);
assign II15999 = ((~g10423))|((~g2683));
assign g6464 = ((~II10398));
assign g10546 = ((~II16203));
assign g6572 = ((~g5805));
assign g7477 = ((~II11869));
assign II6159 = ((~g2123));
assign g9009 = ((~II14405));
assign II15293 = ((~g10001));
assign g10278 = ((~g10182));
assign g8277 = ((~II13203));
assign g5485 = (g1914&g4257);
assign g7913 = ((~g7467));
assign g10717 = (g6235)|(g10705);
assign g2212 = ((~g686));
assign II7920 = ((~g3440));
assign g6048 = ((~II9673));
assign g5531 = (g1666&g4306);
assign g2223 = ((~II5203))|((~II5204));
assign g7144 = ((~II11387));
assign g4670 = (g192&g3946);
assign II9688 = ((~g5201));
assign g8294 = ((~II13236));
assign II16487 = ((~g10771));
assign II5629 = (g845)|(g841)|(g837);
assign II12366 = ((~g7134));
assign g6883 = (g1923&g6413);
assign II11974 = ((~g7001))|((~II11973));
assign g10544 = (g5511)|(g10495);
assign II9338 = ((~g5576));
assign g8890 = ((~II14236));
assign g5035 = ((~II8410));
assign II11296 = ((~g6525));
assign g6803 = ((~II10819));
assign g11021 = (g448&g10974);
assign II6979 = ((~g2888));
assign g11172 = (g486&g11112);
assign g11614 = ((~II17662));
assign g7441 = (g7271)|(g6789);
assign g5524 = (g1678&g4291);
assign g8399 = (g6094&g8229);
assign g10223 = ((~II15595));
assign II8728 = ((~g4605))|((~g1117));
assign II16363 = ((~g10599));
assign g11350 = ((~g11287));
assign g8198 = ((~II13131));
assign g11551 = (g11538&g4013);
assign g10528 = ((~g10464));
assign g8425 = ((~II13589));
assign II13776 = ((~g8513));
assign g9686 = (g9454)|(g9292)|(g9274);
assign II7048 = ((~g2807));
assign g8925 = ((~II14252));
assign g10197 = ((~II15565));
assign II6495 = ((~g2076));
assign II10445 = ((~g5770));
assign II12644 = ((~g7729));
assign g7682 = ((~g7148));
assign g10864 = (g5532)|(g10751);
assign g6655 = (g5296&g5812);
assign II6264 = ((~g2118));
assign g6710 = ((~II10693));
assign g8363 = ((~II13469));
assign g9824 = ((~II14973));
assign g7850 = ((~II12647));
assign g8845 = (g8611&g8711);
assign g7008 = ((~II11149));
assign II9558 = ((~g5598))|((~II9557));
assign II9605 = ((~g5620));
assign g6117 = ((~II9804));
assign II13859 = ((~g1448))|((~II13857));
assign g5166 = ((~g4682));
assign g7388 = ((~II11773));
assign II12229 = ((~g7070));
assign g2024 = ((~g1718));
assign g11219 = (g11145)|(g11006);
assign II7417 = ((~g4160));
assign g4636 = ((~II8036));
assign g7733 = ((~II12380));
assign g11345 = ((~II17158));
assign II12765 = ((~g7638));
assign II5282 = ((~g758))|((~g762));
assign g10751 = (g10646&g4013);
assign g10971 = (g10849&g3161);
assign g7882 = ((~g7479));
assign g8667 = ((~II13952));
assign g6175 = ((~g5320));
assign g8616 = ((~II13868))|((~II13869));
assign g11483 = (g6633)|(g11460);
assign II5728 = ((~g2084));
assign g5821 = ((~II9433));
assign g5143 = ((~g4682));
assign g6930 = (g6364)|(g4269);
assign g5211 = (g1080&g4724);
assign g3052 = ((~II6264));
assign II10274 = ((~g5811));
assign II15214 = (g8170)|(g9906)|(g9935)|(g9831);
assign II6911 = ((~g2825));
assign g10763 = (g10639&g4840);
assign II5926 = ((~g2172));
assign II17312 = ((~g11392));
assign g7317 = ((~II11599));
assign II10282 = ((~g6163));
assign II17306 = ((~g11381))|((~II17305));
assign II11383 = ((~g6385));
assign II12457 = ((~g7559));
assign g5196 = ((~II8605))|((~II8606));
assign g7385 = (g7235)|(g6746);
assign g6085 = ((~II9734));
assign g4467 = ((~g3829));
assign g6720 = ((~II10713));
assign II16000 = ((~g10423))|((~II15999));
assign II8379 = ((~g4231));
assign g9452 = ((~II14645));
assign g10758 = (g10652&g4013);
assign g4805 = ((~g3337));
assign g2273 = ((~g881));
assign II11394 = ((~g6621));
assign g8767 = (g8616&g5151);
assign II14906 = ((~g9508));
assign g6554 = (g5075&g6183);
assign g7849 = ((~II12644));
assign g5245 = ((~g4369));
assign II13314 = ((~g8260));
assign g6450 = ((~II10378));
assign g2917 = (g2424&g1657);
assign g11240 = (g5481&g11111);
assign II11241 = ((~g6760))|((~g790));
assign g110 = ((~II4786));
assign II6487 = ((~g2306))|((~g1227));
assign g2038 = ((~g1776));
assign II13376 = ((~g8226));
assign II13273 = ((~g1918))|((~II13272));
assign g9947 = (g9927&g9392);
assign g5218 = ((~II8647));
assign g6915 = (g6347)|(g5686);
assign g3301 = (g1346&g2544);
assign g4769 = ((~g3586));
assign II14876 = ((~g9526));
assign II14694 = ((~g9259));
assign II7269 = ((~g2851));
assign g7432 = ((~II11824));
assign g10948 = (g2223&g10809);
assign g7331 = ((~II11641));
assign II12376 = ((~g7195));
assign g10771 = (g5533)|(g10684);
assign II15257 = ((~g9984))|((~II15256));
assign g3946 = ((~II7099));
assign g8132 = ((~II12999));
assign g5075 = ((~g4439));
assign g3161 = ((~II6367));
assign II4866 = ((~g579));
assign II16007 = ((~g10424))|((~g2689));
assign g4189 = ((~II7384));
assign II7876 = ((~g4109))|((~II7875));
assign g7357 = ((~II11719));
assign g7965 = ((~II12759));
assign g10126 = ((~II15380));
assign g4093 = ((~g2965));
assign g7188 = ((~II11408));
assign II9046 = ((~g4736));
assign gbuf2 = (g878);
assign g9531 = ((~II14678));
assign II13553 = ((~g668))|((~II13552));
assign II10102 = ((~g5730));
assign g9835 = (g9735&g9785);
assign g10508 = (g10391&g2135);
assign II15162 = ((~g9958));
assign II11614 = ((~g6838));
assign g2407 = ((~g197));
assign g5883 = ((~g5309));
assign g6701 = (g6185&g4228);
assign g2355 = ((~II5435));
assign II7035 = ((~g1868))|((~II7033));
assign II8285 = ((~g4771));
assign g10264 = ((~g10128));
assign g11079 = ((~II16850));
assign II6324 = ((~g1864))|((~II6322));
assign g10779 = ((~II16468))|((~II16469));
assign g8622 = ((~g8485));
assign II7411 = ((~g4140));
assign II5050 = ((~g1216));
assign g1990 = ((~g774));
assign g4789 = ((~g3337));
assign g2646 = ((~g1992));
assign II5469 = ((~g1245))|((~II5468));
assign g7306 = ((~II11566));
assign g8151 = ((~g8036));
assign g2579 = ((~g1969));
assign g2174 = ((~g31));
assign g2542 = ((~g1868));
assign g10454 = (g10435&g3411);
assign II15266 = ((~g10001));
assign II13259 = ((~g1900))|((~II13258));
assign g7342 = ((~II11674));
assign g3729 = ((~II6907));
assign g4436 = ((~g3638));
assign g4509 = ((~II7906));
assign II9096 = ((~g5568));
assign II14579 = ((~g9272));
assign g7269 = ((~II11509))|((~II11510));
assign g5623 = ((~II9053));
assign g10462 = ((~II15977));
assign II11318 = ((~g6488));
assign II13209 = ((~g8198));
assign g11300 = (g11213)|(g11091);
assign II11845 = ((~g6869));
assign II13309 = ((~g617))|((~II13307));
assign g11195 = ((~g11112));
assign g10062 = ((~II15284));
assign II17368 = ((~g11423));
assign g3992 = ((~g2571))|((~g2550))|((~g2990));
assign g11109 = ((~g10974));
assign g7746 = ((~II12403));
assign g3374 = (g1231&g3047);
assign II12442 = ((~g7672));
assign g9928 = (g9870)|(g9717);
assign g4443 = ((~g3359));
assign g3629 = ((~g3228));
assign II6716 = ((~g201))|((~II6714));
assign II8161 = ((~g3637));
assign g4429 = ((~II7779));
assign g10723 = (g4952)|(g10633);
assign II13249 = ((~g1891))|((~II13248));
assign g8814 = (g7945)|(g8728);
assign II13785 = ((~g8516));
assign g5725 = (g1580&g5166);
assign g11296 = (g5482&g11241);
assign II9168 = ((~g5040));
assign g10537 = ((~II16178));
assign g11285 = (g11255)|(g11161);
assign g10141 = ((~II15421));
assign g3586 = (g3323&g2191);
assign g11221 = (g11146)|(g11007);
assign II6569 = ((~g3186));
assign II5932 = ((~g2539));
assign II13089 = ((~g8006))|((~g1840));
assign g3089 = (g2054&g2050);
assign g10091 = ((~II15320));
assign g6622 = (g336&g6165);
assign g6109 = ((~g5052));
assign g10652 = (g10627)|(g7743);
assign II11926 = ((~g6900));
assign g4472 = ((~II7847));
assign II11698 = ((~g7057));
assign II12490 = ((~g7637));
assign g6319 = (g1296&g5949);
assign II7459 = ((~g3720));
assign II16856 = ((~g10909));
assign g3720 = ((~II6888));
assign g11162 = ((~g10950));
assign II11303 = ((~g6526));
assign II17142 = ((~g11301));
assign II7523 = ((~g4095));
assign II5289 = ((~g49));
assign g9877 = ((~g9512)&(~g9536)&(~g9569)&(~II15042));
assign II9256 = ((~g5078));
assign g10153 = ((~II15452))|((~II15453));
assign g9599 = (g8&g9292);
assign g5595 = (g1621&g4524);
assign g8566 = ((~II13791));
assign g8782 = ((~II14083));
assign g3143 = ((~II6363));
assign g10530 = ((~g10466));
assign g9344 = ((~II14537));
assign II5986 = ((~g2194));
assign g3516 = (g1209&g3015);
assign g3458 = ((~g3144));
assign g10148 = ((~g10121));
assign g4053 = (g2701&g2276);
assign II9483 = ((~g5050));
assign II8626 = ((~g511))|((~II8624));
assign II12296 = ((~g7236));
assign II6309 = (g2446&g2451&g2456&g2475);
assign g4975 = ((~II8351));
assign II8903 = ((~g4561));
assign g8921 = (g8827)|(g8748);
assign g11422 = ((~II17321));
assign II5077 = ((~g35));
assign g6940 = (g6472&g1945);
assign II8410 = ((~g4283));
assign g10912 = ((~II16688));
assign II16723 = ((~g10851));
assign g4712 = (g1071&g3638);
assign g4758 = ((~g3586));
assign II8650 = ((~g4824))|((~g778));
assign g11612 = (g11599)|(g11590);
assign II15514 = ((~g10122));
assign g3583 = ((~II6742));
assign g10582 = (g10532&g9473);
assign g6568 = ((~g5797));
assign g6063 = ((~g5446));
assign g8695 = ((~II13978));
assign g7975 = ((~II12773));
assign II9253 = ((~g5052));
assign g6529 = (g5757)|(g5000);
assign g3529 = ((~g2310))|((~g3062))|((~g2325));
assign g6191 = ((~g5446));
assign g10908 = ((~II16676));
assign g5276 = (g736&g4780);
assign II11225 = ((~g6534));
assign II7205 = ((~g2632));
assign g5992 = ((~II9608));
assign g4363 = ((~II7654));
assign g10557 = (g4123)|(g10508);
assign g8077 = ((~II12933));
assign g10376 = ((~g10323)&(~g3113));
assign g9417 = (g1738&g9052);
assign g11093 = (g841&g10950);
assign II14564 = ((~g9026));
assign g6454 = ((~II10388));
assign II16953 = ((~g11082));
assign II12168 = ((~g7256));
assign II9591 = ((~g5095));
assign g7781 = ((~II12508));
assign g8954 = ((~II14315));
assign g4412 = ((~II7746));
assign g11247 = (g11097)|(g10949);
assign g7768 = ((~II12469));
assign g5068 = ((~g4840));
assign g5752 = ((~II9326));
assign g6431 = ((~g6145));
assign g8226 = (g7504)|(g8002);
assign II4995 = ((~g416))|((~g309));
assign g6300 = ((~II10159));
assign g11512 = ((~II17555));
assign II9440 = ((~g5078));
assign II6256 = ((~g2462));
assign II13577 = ((~g8330));
assign II17642 = ((~g11579));
assign g8096 = ((~II12953));
assign II15380 = ((~g10098));
assign g5994 = ((~II9612));
assign g2524 = ((~g986));
assign II13385 = ((~g8230));
assign g10456 = ((~II15959));
assign g4238 = (g3999)|(g4007);
assign II7220 = ((~g3213));
assign g8977 = ((~II14352));
assign II8724 = ((~g4791));
assign II10162 = ((~g5943));
assign g8882 = ((~II14217))|((~II14218));
assign g4417 = ((~II7757));
assign II12196 = ((~g7272));
assign g5696 = ((~II9229));
assign g10353 = ((~II15823));
assign g10137 = ((~II15409));
assign g6558 = ((~II10484));
assign g9151 = (g8967&g6674);
assign g9673 = (g9454)|(g9292)|(g9274);
assign g1999 = ((~g806));
assign II5740 = ((~g2341));
assign II8751 = ((~g4613))|((~II8750));
assign II12849 = ((~g7632));
assign g10905 = ((~II16667));
assign g5823 = (g5631)|(g4882);
assign II5576 = (g431)|(g435)|(g440)|(g444);
assign II15488 = ((~g10116));
assign II12123 = ((~g6861));
assign II12279 = ((~g7225));
assign II17669 = ((~g11604));
assign II11996 = ((~g7107))|((~II11995));
assign g9386 = (g1327&g9151);
assign II5358 = (g1245)|(g1240)|(g1235)|(g1275);
assign II15908 = ((~g10302))|((~II15906));
assign g2549 = ((~g1386));
assign g6398 = ((~II10302));
assign g8357 = ((~II13451));
assign g3354 = (g2920)|(g2124);
assign g6534 = (g5772)|(g5003);
assign II16647 = ((~g10866));
assign g4066 = ((~II7191));
assign g5230 = (g1265&g4735);
assign II10278 = ((~g5815));
assign g8139 = ((~g8025));
assign II6260 = ((~g2025));
assign g4583 = ((~g3880));
assign II7399 = ((~g4113));
assign g6589 = ((~II10549));
assign g4772 = ((~g3440));
assign II9383 = ((~g5296));
assign II15235 = ((~g9968));
assign II16784 = ((~g10895));
assign g10593 = ((~II16264));
assign g4631 = ((~g3820));
assign II10075 = ((~g5724));
assign II11076 = ((~g6649));
assign II9762 = ((~g5276));
assign g7078 = ((~II11309));
assign g3820 = ((~II7048));
assign g8789 = (g8639&g8719);
assign g7903 = ((~g7446));
assign g7043 = ((~II11214));
assign II5149 = ((~g1453));
assign g5476 = (g1615&g4237);
assign g10747 = ((~II16432));
assign II6891 = ((~g2962));
assign II13360 = ((~g8126));
assign g7146 = ((~II11391));
assign g5850 = ((~g5320));
assign II5611 = ((~g1280))|((~g1284));
assign II9208 = ((~g5047));
assign II5843 = ((~g2509));
assign g4366 = ((~II7659));
assign II9087 = ((~g5113));
assign g7096 = (g6544)|(g5911);
assign g7989 = ((~II12805));
assign g10364 = ((~g10327)&(~g3744));
assign g2016 = ((~g1361));
assign g7679 = (g1950&g6863);
assign g7347 = ((~II11689));
assign II11326 = ((~g6660));
assign II13627 = ((~g8326));
assign g6183 = ((~g5320));
assign g9736 = (g9430)|(g9416);
assign II15855 = ((~g10336));
assign II17350 = ((~g11377));
assign g11047 = ((~II16802));
assign g8541 = ((~g4001))|((~g8390));
assign g9527 = ((~II14668));
assign g8445 = ((~II13633));
assign g7010 = ((~II11155));
assign g9509 = (g9151)|(g9125)|(g9111);
assign II17100 = ((~g11221));
assign g4109 = (g806&g3287);
assign g10304 = (g10211&g9079);
assign g4394 = ((~II7729));
assign II11135 = ((~g6679));
assign II13005 = ((~g8046));
assign g10858 = (g5501)|(g10741);
assign g5681 = (g135&g5361);
assign g3275 = (g115&g2356);
assign II14690 = ((~g9150));
assign II9567 = ((~g5556));
assign II6337 = (g201&g2421&g2407&g2396);
assign g6684 = (g5314&g5836);
assign g11332 = (g11273)|(g11172);
assign II13020 = ((~g8049));
assign II17537 = ((~g11497));
assign II13522 = ((~g695))|((~II13521));
assign g11583 = (g1314&g11541);
assign II17636 = ((~g11577));
assign gbuf9 = (g1957);
assign g4292 = ((~g3863));
assign II9479 = ((~g4954));
assign g7312 = ((~II11584));
assign g9866 = (g1549&g9802);
assign g11214 = (g950&g11159);
assign g10627 = (g10548&g4564);
assign II6794 = ((~g143))|((~II6792));
assign II5348 = ((~g746));
assign g8061 = ((~II12901));
assign II9006 = ((~g4492))|((~g1791));
assign II6177 = ((~g2177))|((~II6176));
assign II9013 = ((~g4767));
assign g7609 = ((~II12177));
assign II16087 = ((~g861))|((~II16086));
assign g3268 = (g466&g2511);
assign g7778 = ((~II12499));
assign II6836 = ((~g3287))|((~g806));
assign II11055 = ((~g6419));
assign II13105 = ((~g7929));
assign g3364 = ((~g3121));
assign II17701 = ((~g11617));
assign II5850 = ((~g2273));
assign g5546 = ((~II8973));
assign g6878 = ((~II10966));
assign g5309 = (g3664)|(g4401);
assign II9053 = ((~g4752));
assign II6338 = (g2475&g2456&g2451&g2446);
assign II16149 = (g10472)|(g10470)|(g10468)|(g10467);
assign g7365 = ((~II11743));
assign II17182 = ((~g11309));
assign II5518 = ((~g1019))|((~II5516));
assign II7154 = ((~g2617));
assign g7801 = ((~II12568));
assign g5513 = (g1675&g4282);
assign II13293 = ((~g1882))|((~g8161));
assign g5733 = ((~II9287));
assign g11454 = ((~II17419));
assign g5767 = ((~II9349));
assign g7744 = ((~II12397));
assign g4378 = ((~II7697));
assign II7366 = ((~g4012));
assign II5351 = (g1145)|(g1141)|(g1137)|(g1133);
assign g4340 = (g1153&g3715);
assign g9889 = ((~II15072));
assign g10193 = ((~g10057));
assign g6281 = ((~II10102));
assign g10888 = ((~II16626));
assign g5418 = (g1512&g4344);
assign g7138 = (g6055&g6707);
assign g8309 = ((~II13308))|((~II13309));
assign g10361 = ((~g10268));
assign II12776 = ((~g7586));
assign g2351 = ((~II5427));
assign g8428 = (g8382)|(g8068);
assign g11593 = ((~II17633));
assign g11270 = (g11198)|(g11032);
assign II10153 = ((~g5947));
assign II17228 = ((~g11300));
assign g11005 = (g5119&g10827);
assign II17288 = ((~g11366))|((~g11363));
assign II7342 = ((~g4011));
assign g2228 = ((~g28));
assign g10761 = (g10700&g10699);
assign II8456 = ((~g4472));
assign g3186 = ((~II6373));
assign II9684 = ((~g5426));
assign g10122 = ((~II15374));
assign II16330 = ((~g10616))|((~g4997));
assign g9820 = ((~II14961));
assign g3532 = ((~g3164));
assign g4186 = ((~II7375));
assign g10189 = ((~II15545));
assign g2119 = ((~II5031));
assign g4314 = ((~g4013));
assign g3983 = ((~g3222));
assign g2798 = ((~g2449));
assign g4329 = ((~g4144));
assign g9933 = (g9912&g9624);
assign II11756 = ((~g7191));
assign II17194 = ((~g11317));
assign g9263 = ((~g8892));
assign g7897 = ((~g7712));
assign g4958 = ((~II8328));
assign g7212 = ((~II11444));
assign g3414 = (g2911)|(g2917);
assign g4837 = (g1068&g3638);
assign II6273 = ((~g2482));
assign g10172 = ((~II15510));
assign II16261 = ((~g10556));
assign II15523 = ((~g10058));
assign II5862 = ((~g2537));
assign II4956 = ((~g327))|((~II4954));
assign II15329 = ((~g9995));
assign g4992 = (g1407&g4682);
assign g3406 = ((~II6611));
assign g7359 = ((~II11725));
assign g2853 = ((~g2171));
assign g4004 = ((~II7140));
assign II10651 = ((~g6035));
assign II13828 = ((~g8488));
assign II8715 = ((~g4601))|((~g4052));
assign g8401 = (g677&g8124);
assign g8874 = ((~II14194));
assign g7602 = ((~II12156));
assign II6409 = ((~g2356));
assign g2752 = ((~II5824));
assign g11071 = ((~g10913));
assign g7190 = ((~II11412));
assign II16531 = ((~g10720));
assign g6815 = ((~II10855));
assign g6198 = (g1499&g5128);
assign II9625 = ((~g5405));
assign II17258 = ((~g11345));
assign g9339 = ((~II14522));
assign g7062 = ((~II11262))|((~II11263));
assign II14948 = ((~g9555));
assign g10031 = ((~II15229));
assign II12094 = ((~g1490))|((~II12092));
assign g9713 = (g1589&g9474);
assign g6830 = (g1380&g6596);
assign g8777 = (g5522)|(g8659);
assign g10805 = (g10759)|(g10760);
assign g4380 = ((~II7701));
assign g8747 = ((~II14040));
assign g10144 = ((~II15431))|((~II15432));
assign g6839 = (g1397&g6596);
assign g6228 = (g5605&g713);
assign g9955 = (g9947)|(g9941)|(g9808);
assign g5649 = ((~II9108));
assign II7255 = ((~g3227));
assign g2802 = ((~g2276));
assign g8248 = (g8014)|(g7707);
assign g4551 = ((~g3946));
assign g8821 = (g8643&g8751);
assign g8826 = ((~g8739))|((~g8737))|((~g8648));
assign g4220 = (g105&g3539);
assign g3663 = ((~II6832));
assign II10610 = ((~g5879));
assign g5857 = (g5418)|(g4670);
assign g4488 = ((~II7876))|((~II7877));
assign g8523 = ((~II13732));
assign g8802 = ((~II14127));
assign g10740 = (g10676&g3384);
assign II15503 = ((~g10044));
assign II14202 = ((~g8825))|((~g591));
assign g11181 = ((~II16944));
assign g2421 = ((~g1374));
assign II8133 = ((~g3632));
assign g7197 = ((~II11423));
assign g10869 = ((~II16577));
assign II11873 = ((~g6863));
assign g2118 = ((~g1854));
assign II15601 = ((~g10173));
assign g4951 = ((~II8320));
assign g4456 = ((~g3375));
assign g7670 = ((~II12289));
assign II12363 = ((~g7187));
assign g11058 = (g10933)|(g5280);
assign II8007 = ((~g3829));
assign II11433 = ((~g6424));
assign II11722 = ((~g7034));
assign II6125 = ((~g2215))|((~II6124));
assign g2791 = ((~g2187)&(~g750));
assign II8098 = ((~g3583));
assign g7426 = ((~II11814));
assign g8376 = ((~II13478));
assign II5973 = ((~g2247));
assign g5741 = ((~II9305));
assign II11194 = ((~g6515));
assign II13744 = ((~g8297));
assign g10786 = ((~II16484));
assign g7808 = ((~II12589));
assign g10182 = ((~II15530));
assign II11180 = ((~g6506));
assign g10437 = ((~g10333));
assign g8670 = ((~g8551));
assign g11626 = ((~II17692));
assign g8718 = (g8600&g7903);
assign II7104 = ((~g3186));
assign g7825 = (g1941&g7479);
assign g6913 = ((~II11021));
assign g2432 = ((~II5513));
assign g2268 = ((~g654));
assign II9120 = ((~g5218));
assign g4257 = ((~g3664));
assign II12598 = ((~g7628));
assign g2439 = ((~g1814))|((~g1828));
assign II14400 = ((~g8891));
assign g10724 = (g10312)|(g10672);
assign II12215 = ((~g7061))|((~II12214));
assign g10275 = ((~II15669));
assign g11488 = (g6671)|(g11465);
assign II13816 = ((~g8559));
assign g9310 = ((~II14503));
assign g11601 = (g1351&g11574);
assign g9895 = ((~II15088));
assign II17051 = ((~g10923))|((~g11249));
assign g4371 = ((~II7674));
assign g10414 = (g10300)|(g9534);
assign II7865 = ((~g774))|((~II7863));
assign g4227 = ((~g3292)&(~g3793)&(~g2586)&(~g2579));
assign g4327 = ((~II7600));
assign g9906 = (g9873&g9683);
assign II13122 = ((~g7966));
assign g4536 = ((~g3880));
assign g5391 = ((~II8827));
assign II10769 = ((~g5944))|((~g1801));
assign g5128 = (g4474&g2733);
assign g4749 = ((~g3710))|((~g2061));
assign II14211 = ((~g599))|((~II14209));
assign g4335 = ((~II7612));
assign g6618 = (g658&g6016);
assign II7450 = ((~g3704));
assign g9091 = ((~g8892));
assign II16534 = ((~g10747));
assign II5258 = ((~g67));
assign g8945 = (g8801)|(g8710);
assign g4195 = ((~II7402));
assign g8764 = (g7443&g8684);
assign II13077 = ((~g1872))|((~II13076));
assign g2275 = ((~g757));
assign g6729 = ((~II10724));
assign g7354 = ((~II11710));
assign g8562 = ((~II13779));
assign g5910 = (g5023)|(g4341);
assign g8240 = ((~g7972));
assign g9422 = (g1750&g9030);
assign g2818 = ((~II5922));
assign II8199 = ((~g4013));
assign II4873 = ((~g105));
assign g6321 = (g1284&g5949);
assign g2813 = ((~II5913));
assign g5222 = ((~g4640));
assign g5233 = (g1791&g4492);
assign g3273 = ((~II6448))|((~II6449));
assign II10771 = ((~g1801))|((~II10769));
assign g6206 = (g560&g5068);
assign g10428 = ((~g10335)&(~g4620));
assign II15986 = ((~g10417));
assign II12004 = ((~g153))|((~II12002));
assign g8449 = ((~II13645));
assign II11289 = ((~g6508));
assign II15284 = ((~g10034));
assign II16370 = ((~g10592));
assign g7546 = ((~II11970));
assign II12910 = ((~g7922));
assign g3522 = ((~g3164));
assign II13099 = ((~g7927));
assign II13902 = ((~g1428))|((~II13900));
assign II7662 = ((~g3336));
assign g7001 = ((~II11140));
assign g10050 = ((~II15269));
assign g5001 = (g1300&g4491);
assign g5171 = ((~II8562))|((~II8563));
assign II13894 = ((~g8529))|((~II13893));
assign II11357 = ((~g6594));
assign g9108 = ((~II14449));
assign g3989 = (g248&g3164);
assign g7633 = ((~II12239));
assign g3434 = (g237&g3228);
assign g3710 = ((~g3215));
assign g3256 = ((~II6424));
assign g2908 = ((~II6077));
assign II8762 = ((~g4616))|((~II8761));
assign II12829 = ((~g7680));
assign II6421 = ((~g2346));
assign g8797 = ((~II14116));
assign g10263 = ((~g10127));
assign g5703 = (g174&g5361);
assign II17695 = ((~g11614));
assign g7067 = ((~II11279))|((~II11280));
assign g8639 = (g8118)|(g8462);
assign g8066 = ((~II12916));
assign g4006 = (g201&g3228);
assign II16769 = ((~g10894));
assign II6436 = ((~g2351));
assign g8576 = ((~II13819));
assign g5642 = ((~II9087));
assign g2892 = (g1980&g1976);
assign g5848 = (g3860&g5519);
assign g7815 = ((~II12610));
assign g2096 = ((~II4929))|((~II4930));
assign g11628 = ((~II17698));
assign II7713 = ((~g3750));
assign g2743 = ((~II5801));
assign II15708 = ((~g10241));
assign g10252 = ((~g10137));
assign g10281 = ((~g10162));
assign g2166 = ((~II5101));
assign g4430 = ((~II7782));
assign II13185 = ((~g8192));
assign g8783 = ((~g8746));
assign II14552 = ((~g9264));
assign g8984 = ((~II14373));
assign g1981 = ((~g650));
assign g11656 = ((~II17770));
assign g8047 = (g7557&g5919);
assign g2073 = ((~II4879));
assign g7628 = ((~II12226));
assign II17487 = ((~g11474))|((~II17485));
assign II8192 = ((~g3566));
assign g6313 = ((~II10198));
assign II17268 = ((~g11351));
assign g8711 = ((~g8677));
assign II17295 = ((~g11373))|((~g11369));
assign g5836 = ((~g5320));
assign g11445 = ((~II17384));
assign II16059 = ((~g841))|((~II16058));
assign II5323 = ((~g1336))|((~g1341));
assign II6553 = ((~g3186));
assign g4763 = ((~g3586));
assign II17321 = ((~g11348));
assign g10203 = ((~g10177));
assign II17681 = ((~g11608));
assign II17401 = ((~g11418))|((~II17400));
assign g4500 = (g1357&g3941);
assign g8628 = ((~II13894))|((~II13895));
assign g9859 = (g9736&g9573);
assign g6956 = ((~II11106));
assign g7224 = (g5398&g6441);
assign g11407 = (g11339&g5949);
assign II14303 = ((~g8811));
assign g9870 = (g1561&g9816);
assign g7753 = ((~II12424));
assign II11508 = ((~g6580))|((~g1806));
assign II11501 = ((~g6581));
assign g6751 = ((~II10762));
assign II16379 = ((~g10598));
assign g6240 = (g182&g5361);
assign g10297 = (g8892&g10211);
assign g5529 = (g4129&g4288);
assign II9662 = ((~g5319));
assign II17188 = ((~g11313));
assign g6693 = (g5494&g5845);
assign II12003 = ((~g7082))|((~II12002));
assign g9651 = (g944&g9240);
assign II9248 = ((~g4954));
assign g3261 = ((~g2229))|((~g2222))|((~g2211))|((~g2202));
assign II7185 = ((~g2626));
assign g4609 = (g3400)|(g119);
assign g8415 = ((~II13560))|((~II13561));
assign g8598 = (g8471&g7432);
assign g8162 = (g7898)|(g6889);
assign II13329 = ((~g8116));
assign g3815 = ((~g3228));
assign II6576 = ((~g2617));
assign g10307 = ((~II15729));
assign g2555 = ((~II5676))|((~II5677));
assign II7233 = ((~g2817));
assign g6842 = ((~II10898));
assign g8602 = (g8401)|(g8550);
assign g10430 = ((~g10349)&(~g3566));
assign g4205 = ((~II7432));
assign II13367 = ((~g8221));
assign II10813 = ((~g6397));
assign g4561 = (g538&g4003);
assign g6514 = (g5738)|(g4992);
assign g5201 = (g1250&g4721);
assign g6151 = ((~II9872));
assign g4558 = ((~g3880));
assign g3756 = ((~g3015));
assign g6361 = ((~g5867));
assign g11103 = (g2250&g10937);
assign II7276 = ((~g2861));
assign g6644 = ((~II10601));
assign II10901 = ((~g6620));
assign II10394 = ((~g5824));
assign g7071 = (g5916&g6590);
assign g7200 = (g3098&g6418);
assign g2001 = ((~g814));
assign g4949 = (g3505&g4449);
assign g10393 = ((~g10317));
assign II13347 = ((~g8122));
assign g11387 = (g11284&g3629);
assign g8342 = ((~II13406));
assign g9775 = ((~g9474));
assign II12655 = ((~g7402));
assign II8985 = ((~g4733));
assign g6705 = ((~II10682));
assign g7998 = ((~II12822));
assign g5193 = ((~g4682));
assign g1973 = ((~g466));
assign g10347 = ((~II15807));
assign g8790 = ((~II14101));
assign g2084 = ((~II4900));
assign g4783 = ((~g3829));
assign II13338 = ((~g8210));
assign g11390 = ((~II17219));
assign g2777 = ((~g2276));
assign g5575 = (g1618&g4501);
assign II9810 = ((~g5576));
assign g10521 = (II16148)|(II16149);
assign II12517 = ((~g7737));
assign g4492 = (g1786&g3685);
assign g6014 = ((~g5309));
assign g5892 = ((~II9519));
assign g2296 = ((~II5332));
assign II5341 = ((~g315))|((~g426));
assign g4306 = ((~g3586));
assign II14140 = ((~g8717));
assign II13513 = ((~g686))|((~g8248));
assign II13388 = ((~g8230));
assign g7723 = ((~II12354));
assign II8604 = ((~g4259))|((~g506));
assign g7327 = ((~II11629));
assign g4575 = ((~g3880));
assign II7213 = ((~g2635));
assign g9649 = (g916&g9205);
assign II9368 = ((~g5288));
assign g7039 = ((~II11204));
assign g4889 = ((~II8240));
assign g11050 = ((~II16811));
assign g4512 = (g357&g3586);
assign II10719 = ((~g6003));
assign g10576 = ((~g10524));
assign g8175 = (g5291&g7853);
assign II8293 = ((~g4779));
assign II13878 = ((~g1444))|((~II13876));
assign g6715 = ((~II10702));
assign g7205 = ((~II11433));
assign g9841 = (g9706&g9512);
assign II14277 = ((~g8847))|((~g1828));
assign II13166 = ((~g8009));
assign g5052 = ((~g4394));
assign II17413 = ((~g11425));
assign g4010 = ((~g3144));
assign II8204 = ((~g3976));
assign g4896 = ((~II8253));
assign g8510 = (g8414&g7972);
assign II9901 = ((~g5557));
assign g5612 = (g1627&g4543);
assign g2013 = ((~g1101));
assign g5444 = (g1041&g4880);
assign II9930 = ((~g5317));
assign g10250 = ((~g10136));
assign II16811 = ((~g10908));
assign g5148 = (g3088&g4671);
assign g7587 = ((~II12086))|((~II12087));
assign g4874 = ((~II8215));
assign g7520 = ((~II11898));
assign g9585 = (g889&g8995);
assign II12571 = ((~g7509));
assign g5280 = (g4593&g3052);
assign II5279 = ((~g73));
assign g5179 = ((~II8576))|((~II8577));
assign II7249 = ((~g2833));
assign g6299 = ((~II10156));
assign II13711 = ((~g8342));
assign g8800 = ((~II14123));
assign g10464 = ((~II15983));
assign II6666 = ((~g2776))|((~II6664));
assign II12403 = ((~g7611));
assign g10408 = (g10298)|(g9553);
assign g2593 = ((~g1973));
assign g8677 = ((~II13962));
assign g3212 = ((~II6385));
assign II10072 = ((~g5719));
assign g11299 = (g5498&g11243);
assign II10381 = ((~g5847));
assign g6258 = ((~II10033));
assign g10895 = ((~II16647));
assign g8427 = ((~II13595));
assign II15171 = (g8175)|(g9909)|(g9896)|(g9835);
assign g3215 = ((~g2564))|((~g1822));
assign II12484 = ((~g7580));
assign II11173 = ((~g6500));
assign II17510 = ((~g11481));
assign g5737 = (g1524&g5183);
assign g5812 = ((~g5320));
assign II7447 = ((~g3694));
assign g3208 = ((~II6381));
assign g6262 = ((~II10045));
assign g3681 = ((~II6837))|((~II6838));
assign g4882 = (g1089&g3638);
assign g6231 = (g818&g5608);
assign g3914 = ((~g3015));
assign II17742 = ((~g11636));
assign g2330 = ((~g1891));
assign II10221 = ((~g6117));
assign g6123 = (g5630&g4311);
assign II5245 = ((~g925));
assign g6592 = (g5100)|(g5882);
assign g10494 = (g10433&g3945);
assign g6336 = ((~II10231));
assign g6171 = ((~g5446));
assign g8213 = ((~g7826));
assign II5497 = ((~g587));
assign g7534 = ((~II11942));
assign g10233 = ((~g10187));
assign g7263 = ((~II11498));
assign g10268 = (g10183&g3307);
assign g6798 = ((~II10804));
assign II16046 = ((~g10370))|((~II16044));
assign II11731 = ((~g7021));
assign II17749 = ((~g11644));
assign g8965 = (g8110&g6778&g8849);
assign g9915 = (g9853)|(g9693);
assign g9367 = (g9335)|(g9331);
assign II9265 = ((~g5085));
assign g11632 = ((~II17710));
assign II10138 = ((~g5677));
assign g10791 = (g6186)|(g10762);
assign g6901 = (g6788)|(g6247);
assign g2728 = ((~g2025));
assign g2057 = ((~g754));
assign g3105 = ((~g2482));
assign II10084 = ((~g5742));
assign II9801 = ((~g5416));
assign II12012 = ((~g6916));
assign g10377 = ((~II15855));
assign g2086 = ((~II4906));
assign g5050 = ((~II8429));
assign g11038 = ((~II16775));
assign g5184 = ((~g4682));
assign g5794 = ((~II9394));
assign g9290 = ((~II14494));
assign g3861 = ((~II7054));
assign g11538 = ((~II17568))|((~II17569));
assign g11509 = ((~II17546));
assign g7296 = (g7131)|(g6322);
assign g4128 = (g1976&g2779);
assign g3939 = (g213&g3164);
assign g8699 = (g7595&g8579);
assign g6746 = (g6228&g6166);
assign II4980 = ((~g333))|((~II4978));
assign g2981 = (g1776&g2264);
assign g5304 = ((~II8779))|((~II8780));
assign II14802 = ((~g9666));
assign II10526 = ((~g6161));
assign g10214 = ((~II15586));
assign g4117 = ((~g3041))|((~g3061));
assign g6107 = ((~II9776));
assign g8381 = ((~II13489));
assign g8023 = (g7367&g7430);
assign g2775 = ((~II5862));
assign g8486 = ((~g8348));
assign II9185 = ((~g4915));
assign II17466 = ((~g11447));
assign g11500 = ((~II17519));
assign g7794 = ((~II12547));
assign g7235 = (g6663&g6447);
assign g6158 = ((~II9883));
assign g9737 = (g9657)|(g9658)|(g9655);
assign g11160 = ((~g10950));
assign g9843 = (g9711&g9519);
assign g4759 = (g406&g3392);
assign II17569 = ((~g1610))|((~II17567));
assign g6330 = ((~II10221));
assign g4714 = (g646&g3333);
assign II9727 = ((~g5250));
assign II13765 = ((~g731))|((~g8417));
assign g6295 = ((~II10144));
assign g2650 = ((~g2006));
assign g8124 = ((~g8011));
assign g4677 = ((~g3501)&(~g2669)&(~g3485)&(~g2655));
assign g6974 = ((~g6365));
assign g9273 = ((~II14490));
assign g3384 = ((~g3143));
assign II8820 = ((~g4473));
assign g7664 = (g6855)|(g4084);
assign II8563 = ((~g491))|((~II8561));
assign g11267 = (g11192)|(g11029);
assign g8055 = (g7588&g5128);
assign II16598 = ((~g10804));
assign g4169 = (g2765&g3066);
assign g6312 = ((~II10195));
assign II13735 = ((~g8293));
assign II6046 = ((~g2218));
assign II10174 = ((~g5994));
assign g9980 = ((~II15181));
assign II8740 = ((~g1121))|((~II8738));
assign g8280 = ((~II13212));
assign g9863 = (g9740&g9576);
assign g10135 = ((~II15403));
assign g11330 = (g11304)|(g11170);
assign II13915 = ((~g8451));
assign g10238 = ((~g10191));
assign g4059 = (g1756&g2796);
assign g4752 = (g401&g3385);
assign g8937 = (g8786)|(g8698);
assign g2695 = ((~g2039));
assign II16982 = ((~g11088));
assign g8019 = (g7386&g4332);
assign g11572 = ((~g11561));
assign II15580 = ((~g10155));
assign g4277 = ((~g3688));
assign g10295 = (g8892&g10208);
assign II14490 = ((~g8885));
assign g4548 = (g440&g3990);
assign II16475 = ((~g10765));
assign g2320 = ((~g18));
assign II12258 = ((~g7103));
assign g8756 = (g7431&g8674);
assign g3630 = ((~II6789));
assign g2003 = ((~g822));
assign II9720 = ((~g5248));
assign II11097 = ((~g6748));
assign g8107 = (g6226&g7882);
assign g9777 = ((~g9474));
assign II13260 = ((~g8153))|((~II13258));
assign II12068 = ((~g7116))|((~II12067));
assign II10180 = ((~g6107));
assign II5638 = ((~g936));
assign II11367 = ((~g6392));
assign g10708 = ((~II16387));
assign g5656 = ((~II9129));
assign g8316 = ((~II13332));
assign g5667 = ((~II9162));
assign g6892 = (g6472&g5805);
assign II14751 = (g8995)|(g9205)|(g9192);
assign g3770 = ((~II6985));
assign g5102 = ((~II8476));
assign g8142 = ((~II13023));
assign g11461 = (g11429&g5446);
assign g8000 = ((~g7011))|((~g7574))|((~g7562))|((~g7550));
assign g5265 = ((~g4362));
assign g7613 = (g6940&g5984);
assign II5023 = ((~g995))|((~g1275));
assign g9705 = (g1580&g9474);
assign II15820 = ((~g10204));
assign g7338 = ((~II11662));
assign II5316 = ((~g1032))|((~II5315));
assign II11068 = ((~g6426));
assign g11233 = (g11085)|(g10946);
assign g2496 = (g374&g369);
assign g3512 = (g2050&g2971);
assign II8892 = ((~g4554));
assign g7241 = (g6772&g6172);
assign g10502 = (g4169)|(g10365);
assign II15725 = ((~g10251));
assign II9068 = ((~g4768));
assign g9904 = (g9886&g9676);
assign II5719 = ((~g2072));
assign g3539 = ((~g3015));
assign II5057 = ((~g1961));
assign g4386 = ((~II7713));
assign g5292 = ((~g4445));
assign g2178 = ((~g45));
assign g6115 = ((~II9798));
assign II6363 = ((~g2459));
assign II8842 = ((~g4556));
assign II10234 = ((~g6114));
assign II12817 = ((~g7692));
assign g4477 = (g1129&g3878);
assign g4373 = ((~II7680));
assign II12796 = ((~g7543));
assign g4552 = ((~g3880));
assign II17161 = ((~g11314));
assign g7427 = ((~II11817));
assign g11017 = ((~II16742));
assign g9833 = (g9729&g9785);
assign g2955 = ((~II6156));
assign II11387 = ((~g6672));
assign g5724 = ((~II9268));
assign g4736 = (g396&g3379);
assign II13280 = ((~g8250));
assign II9749 = ((~g5266));
assign g6795 = (g5036&g5878);
assign g11257 = (g11234)|(g11019);
assign II12107 = ((~g7113))|((~II12106));
assign g8517 = ((~II13720));
assign g7879 = (g7610&g3798);
assign II5449 = ((~g1235))|((~g991));
assign g6277 = ((~II10090));
assign II10126 = ((~g5682));
assign g11010 = (g5187&g10827);
assign II12047 = ((~g1486))|((~II12045));
assign II6523 = ((~g2819));
assign II6168 = ((~g153))|((~II6166));
assign g7410 = ((~II11790));
assign II11494 = ((~g6574));
assign II4900 = ((~g583));
assign II5092 = ((~g32));
assign II13857 = ((~g8538))|((~g1448));
assign g10259 = ((~g10141));
assign g2944 = (g2424&g1669);
assign g10738 = (g10692&g4840);
assign II6449 = ((~g1776))|((~II6447));
assign g6100 = ((~II9759));
assign g11645 = ((~II17739));
assign g10329 = ((~II15775));
assign g6810 = ((~II10840));
assign g2410 = ((~g1453));
assign g5518 = (g4317&g3532);
assign g4337 = ((~g4144));
assign II6351 = (g2405)|(g2389)|(g2380)|(g2372);
assign g5773 = ((~II9359));
assign II11683 = ((~g7069));
assign g2105 = ((~II4972))|((~II4973));
assign II15453 = ((~g10051))|((~II15451));
assign g8122 = ((~II12981));
assign g8129 = ((~g8015));
assign II15826 = ((~g10205));
assign g6110 = ((~II9783));
assign g6993 = ((~II11135));
assign g8509 = ((~g8366));
assign g6352 = (g278&g5894);
assign II10930 = ((~g6395))|((~g5555));
assign g10927 = ((~g10827));
assign g2172 = ((~g43));
assign g2689 = ((~g2038));
assign II12712 = ((~g7441));
assign g3390 = ((~g3161));
assign II9452 = ((~g5085));
assign g11271 = (g5624&g11191);
assign II10087 = ((~g5753));
assign II14412 = ((~g8939));
assign g8644 = (g8123)|(g8464);
assign II4930 = ((~g321))|((~II4928));
assign g9624 = (g9316)|(g9313);
assign II13945 = ((~g8488));
assign II15872 = ((~g2713))|((~II15870));
assign g8943 = (g8837)|(g8749);
assign g5226 = ((~II8670))|((~II8671));
assign g6506 = (g5731)|(g4989);
assign g11410 = ((~II17271));
assign g7847 = ((~II12638));
assign II13621 = ((~g8315));
assign g7712 = (g7125)|(g3540);
assign g4211 = ((~II7450));
assign g2156 = ((~II5073));
assign g3369 = ((~II6557));
assign II8929 = ((~g4582));
assign II5798 = ((~g2085));
assign II11759 = ((~g7244));
assign g6699 = (g6177&g4221);
assign II5486 = ((~g1011))|((~II5484));
assign g9837 = (g9697&g9751);
assign g8931 = (g8807&g8164);
assign g4158 = ((~g3304));
assign g7284 = ((~II11528));
assign II11914 = ((~g6935))|((~g1494));
assign II5946 = ((~g2176));
assign g10155 = ((~II15461));
assign II9536 = ((~g5008));
assign g4080 = ((~g2903));
assign II16015 = ((~g10425))|((~g2695));
assign II10914 = ((~g6728));
assign g9420 = (g1747&g9030);
assign g2271 = ((~g877));
assign g9272 = (g8934&g3424);
assign g6181 = ((~g5426));
assign g7304 = ((~II11560));
assign g4308 = ((~g3863));
assign II15392 = ((~g10104));
assign g5638 = ((~II9077));
assign g3750 = ((~II6941));
assign II7014 = ((~g2919));
assign II6417 = ((~g2344));
assign g7186 = (g2503&g6403);
assign g6925 = ((~II11043));
assign g2123 = ((~II5047));
assign II17394 = ((~g11415))|((~II17393));
assign g6446 = ((~II10370));
assign g10662 = (g8892&g10571);
assign II11510 = ((~g1806))|((~II11508));
assign g4445 = ((~II7803));
assign g10849 = ((~g10739)&(~g3903));
assign g2207 = ((~II5174));
assign g11040 = ((~II16781));
assign g9328 = (g8971&g5708);
assign g10510 = (g10393&g2135);
assign g1968 = ((~g369));
assign II15247 = ((~g10032));
assign g5533 = (g1724&g4308);
assign II10063 = ((~g5766));
assign g5604 = ((~II9032));
assign II13660 = ((~g1945))|((~II13659));
assign g8332 = ((~II13376));
assign II12607 = ((~g7633));
assign II9866 = ((~g5274));
assign II10864 = ((~g6634));
assign g6075 = (g549&g5613);
assign II7323 = ((~g1231))|((~II7321));
assign g2867 = ((~II6007));
assign g3336 = ((~II6523));
assign II10852 = ((~g6751));
assign II6856 = ((~g3318));
assign II6999 = ((~g2905));
assign g6730 = (g1872&g6128);
assign g6307 = ((~II10180));
assign g7963 = (g7687)|(g7182);
assign g5881 = ((~g5361));
assign g8796 = (g8645&g8725);
assign g9946 = (g9926&g9392);
assign g5895 = ((~g5361));
assign g11068 = ((~g10974));
assign II16635 = ((~g10862));
assign g2445 = ((~II5539))|((~II5540));
assign g3497 = (g2804&g1900);
assign g6253 = ((~II10018));
assign II5292 = ((~g76));
assign g3904 = (g2948&g2779);
assign II11299 = ((~g6727));
assign II16688 = ((~g10800));
assign II14264 = ((~g8843))|((~II14263));
assign g8304 = ((~II13280));
assign II13552 = ((~g668))|((~g8262));
assign g9612 = (g2652&g9240);
assign g5108 = (g1801&g4614);
assign g11615 = (g11601)|(g11592);
assign g4915 = ((~g4413));
assign g2190 = ((~II5149));
assign g7511 = (g6890)|(g6438);
assign g10721 = (g10306)|(g10669);
assign II5020 = ((~g1176));
assign II16616 = ((~g10796));
assign II6489 = ((~g1227))|((~II6487));
assign g2889 = ((~II6049));
assign g10506 = (g10390&g2135);
assign g2827 = ((~g2164));
assign g8431 = (g8387)|(g8071);
assign g5011 = ((~II8385));
assign g6821 = (g237&g6596);
assign g11007 = (g5147&g10827);
assign g4679 = ((~g4013));
assign II8126 = ((~g3662));
assign g8564 = ((~II13785));
assign II6474 = ((~g2297));
assign g11298 = (g11212)|(g11087);
assign g8134 = ((~II13005));
assign g8648 = (g4588&g8511);
assign II12475 = ((~g7545));
assign g3784 = ((~g2586));
assign II13302 = ((~g8162))|((~II13300));
assign II16067 = ((~g2765))|((~II16065));
assign g3734 = ((~g3039))|((~g599));
assign g3141 = ((~g2563));
assign II5371 = ((~g971))|((~g976));
assign g6742 = ((~g5830));
assign g6876 = (g4070&g6560);
assign g5889 = ((~II9514));
assign II11581 = ((~g6826));
assign g5345 = ((~g2754)&(~g4835));
assign g4364 = (g1215&g3756);
assign II13717 = ((~g8354));
assign g4427 = ((~g3638));
assign II10499 = ((~g6149));
assign g6898 = (g6790)|(g4881);
assign g6441 = ((~g6151));
assign g6481 = (g5722)|(g4972);
assign g9875 = ((~II15036));
assign II11065 = ((~g6750));
assign g9392 = (g9328)|(g9324);
assign II5675 = ((~g1218))|((~g1223));
assign g10044 = ((~II15263));
assign g5662 = ((~II9147));
assign g6703 = ((~II10678));
assign II11423 = ((~g6488));
assign II12853 = ((~g7638));
assign g4470 = ((~II7843));
assign g4973 = (g1645&g4467);
assign g2254 = ((~g131));
assign g6620 = ((~II10573));
assign g11077 = ((~g10970)&(~g10971));
assign II17492 = ((~g11475))|((~g3623));
assign g11499 = ((~II17516));
assign II13546 = ((~g8259))|((~II13544));
assign g3732 = ((~II6914));
assign g3944 = ((~g2920));
assign g7454 = ((~g7148));
assign II14097 = ((~g8773));
assign g8951 = ((~II14306));
assign g7951 = (g2868&g7505);
assign g5259 = (g627&g4739);
assign g2855 = ((~II5989));
assign II9642 = ((~g5229));
assign g4264 = (g4048)|(g4053);
assign II11408 = ((~g6405));
assign g11193 = ((~g11112));
assign g4779 = (g501&g3427);
assign II6299 = ((~g2242));
assign g4507 = ((~g3546));
assign II6507 = ((~g2808));
assign g2214 = ((~g115));
assign g7941 = ((~g7406));
assign II13036 = ((~g8053));
assign g10853 = ((~g10731))|((~g5034));
assign g9419 = (g1744&g9030);
assign g8654 = (g8529&g4013);
assign g6885 = ((~II10979));
assign g5066 = ((~II8436));
assign g10166 = ((~II15494));
assign g6405 = ((~g6133));
assign g5746 = (g1589&g5193);
assign g11544 = (g11515&g10584);
assign g2884 = ((~II6040));
assign g10001 = (II15204)|(II15205);
assign g7885 = (g7614&g3812);
assign II17460 = ((~g11449))|((~II17459));
assign g10598 = ((~II16273));
assign II10484 = ((~g6155));
assign g6634 = ((~II10589));
assign II9293 = ((~g5486));
assign II11833 = ((~g7077));
assign II12562 = ((~g7377));
assign g7142 = ((~II11383));
assign g2050 = ((~g1861));
assign g2221 = ((~II5198));
assign g4731 = ((~II8085));
assign g10385 = ((~g10321)&(~g2998));
assign g2044 = ((~II4850));
assign II11531 = ((~g7126));
assign II15424 = ((~g10080));
assign II9080 = ((~g4775));
assign II12948 = ((~g8019));
assign g6083 = (g552&g5619);
assign II11659 = ((~g7097));
assign g6346 = (g5038&g5883);
assign II17549 = ((~g11501));
assign g4616 = ((~g3077)&(~g3491)&(~g2662)&(~g3479));
assign II8480 = ((~g4455))|((~II8479));
assign II13797 = ((~g8473));
assign g10548 = ((~II16209));
assign II17096 = ((~g11219));
assign g2241 = ((~g722));
assign g5504 = ((~g4419));
assign g4725 = (g1032&g3914);
assign II11127 = ((~g6452));
assign g7102 = (g6550)|(g5915);
assign II8328 = ((~g4801));
assign g5627 = ((~g4840));
assign g3584 = (g2863)|(g2516);
assign II4997 = ((~g309))|((~II4995));
assign II11947 = ((~g6905));
assign II16763 = ((~g10890));
assign II7749 = ((~g3764));
assign g8923 = (g8846)|(g8763);
assign II17459 = ((~g11449))|((~g11448));
assign g7766 = ((~II12463));
assign g6286 = ((~II10117));
assign g7048 = ((~II11225));
assign II7033 = ((~g3089))|((~g1868));
assign g10107 = ((~II15341));
assign g8502 = ((~g2382))|((~g605))|((~g591))|((~g8366));
assign g11170 = (g525&g11112);
assign g5030 = (g1280&g4523);
assign II10334 = ((~g6003));
assign g7984 = ((~II12796));
assign g11402 = ((~II17249));
assign II11235 = ((~g6538));
assign g5261 = ((~g4640));
assign g2204 = (g1393)|(g1394);
assign g7755 = ((~II12430));
assign g10331 = (g10256&g3307);
assign II16098 = ((~g10369));
assign II15768 = ((~g10249));
assign g6656 = (g2733&g6061&g4631);
assign g3417 = ((~II6624));
assign g10866 = (g5539)|(g10753);
assign g8380 = (g8252&g4240);
assign g10777 = (g10733&g3015);
assign g4282 = ((~g4013));
assign g10604 = ((~II16280));
assign g9740 = (g9418)|(g9505);
assign g4194 = ((~II7399));
assign g4510 = ((~II7909));
assign g4823 = (g207&g3946);
assign g5865 = ((~II9486));
assign II6879 = ((~g3301))|((~g1351));
assign II5007 = ((~g312))|((~II5005));
assign II5395 = ((~g892));
assign g7363 = ((~II11737));
assign g7731 = ((~II12376));
assign II17522 = ((~g11485));
assign g7956 = ((~g7432));
assign g4140 = ((~II7284));
assign g9807 = ((~g9490));
assign g11020 = (g452&g10974);
assign g5111 = ((~II8499));
assign g8582 = ((~II13825));
assign g11369 = ((~II17194));
assign g3335 = ((~II6520));
assign g3092 = ((~g2181));
assign II14312 = ((~g8814));
assign II15598 = ((~g10170));
assign g6224 = (g1520&g5151);
assign g6980 = ((~II11127));
assign g10526 = ((~g10460));
assign g4284 = ((~g3664));
assign II8835 = ((~g4791));
assign II14379 = ((~g8961));
assign g7460 = ((~g7148));
assign g5819 = (g5625)|(g4876);
assign II9854 = ((~g5557));
assign II6322 = ((~g2050))|((~g1864));
assign g6462 = ((~II10394));
assign II10716 = ((~g6093));
assign g8059 = (g7592&g5919);
assign II16469 = ((~g10518))|((~II16467));
assign g7439 = ((~II11833));
assign II11783 = ((~g7246));
assign g2068 = ((~II4866));
assign g8660 = ((~II13945));
assign g7467 = ((~g7148));
assign II7674 = ((~g3352));
assign g5098 = ((~g4840));
assign g3875 = (g3275)|(g12);
assign II10601 = ((~g5996));
assign g11360 = ((~II17185));
assign g3352 = ((~II6538));
assign II10713 = ((~g6003));
assign g7345 = ((~II11683));
assign II17296 = ((~g11373))|((~II17295));
assign II8215 = ((~g3981));
assign g8255 = ((~g7986));
assign g8365 = (g668&g8240);
assign g6082 = ((~II9727));
assign II15464 = ((~g10094));
assign II10340 = ((~g6205));
assign g6672 = (g5941)|(g5259);
assign g11261 = (g11238)|(g11023);
assign II13674 = ((~g8304));
assign g6089 = ((~g4977));
assign g6967 = ((~II11119));
assign g6777 = (g5691)|(g5052);
assign g9030 = (g8935&g7192);
assign g5037 = ((~II8414));
assign II12303 = ((~g7242));
assign g7915 = ((~g7473));
assign II6034 = ((~g2210));
assign II9896 = ((~g5295));
assign g7472 = (g7148&g2829);
assign g8224 = (g1882&g7887);
assign II8934 = ((~g4271));
assign II12835 = ((~g7660));
assign g7708 = ((~II12339));
assign g6960 = ((~II11112));
assign g2950 = (g2424&g1666);
assign g11095 = (g845&g10950);
assign g2759 = ((~II5843));
assign g4738 = ((~g3440));
assign g4338 = (g1157&g3707);
assign g8611 = (g8410)|(g8556);
assign g3706 = (g471&g3268);
assign II9029 = ((~g4781));
assign g11327 = (g11297)|(g11167);
assign g8196 = ((~II13125));
assign II13433 = ((~g8181));
assign g3759 = ((~II6958));
assign g10370 = ((~g10343)&(~g3463));
assign g11639 = (g11612&g7897);
assign g10355 = ((~II15829));
assign g9343 = ((~II14534));
assign II7654 = ((~g3728));
assign II7099 = ((~g3228));
assign g2374 = ((~g591));
assign g7684 = ((~g7148));
assign g3056 = ((~g2374))|((~g599));
assign g7020 = ((~II11159));
assign II12586 = ((~g7561));
assign g2444 = ((~g876));
assign g7288 = ((~II11540));
assign g8063 = ((~II12907));
assign g9414 = (g1730&g9052);
assign g10807 = (g10701)|(g10761);
assign II13708 = ((~g8337));
assign g10226 = ((~II15598));
assign II13779 = ((~g8514));
assign g11508 = ((~II17543));
assign g2095 = ((~g143));
assign II6838 = ((~g806))|((~II6836));
assign g8273 = ((~II13191));
assign g7509 = ((~II11889));
assign II4859 = ((~g578));
assign II8403 = ((~g4264));
assign g4324 = ((~g4144));
assign g6712 = ((~g5984));
assign g3322 = ((~II6488))|((~II6489));
assign II11989 = ((~g6919));
assign II12978 = ((~g8040));
assign II6757 = ((~g2732));
assign g2185 = ((~g46));
assign g9829 = (g9723&g9785);
assign g6686 = ((~II10651));
assign II11710 = ((~g7020));
assign g6471 = (g5224&g6014);
assign II14982 = ((~g9672));
assign g11334 = (g11277)|(g11174);
assign II9848 = ((~g5557));
assign g8253 = (g8023)|(g7718);
assign II5919 = ((~g2530));
assign g11381 = ((~II17206));
assign g4397 = (g3475&g2181);
assign II15386 = ((~g10101));
assign g2920 = ((~g2462));
assign II17567 = ((~g11496))|((~g1610));
assign II8803 = ((~g4677))|((~g1113));
assign II11444 = ((~g6653));
assign g9529 = ((~II14672));
assign g10868 = ((~II16574));
assign II6770 = ((~g3257))|((~g382));
assign g7360 = ((~II11728));
assign g8049 = (g7567&g5919);
assign g4944 = ((~g4430));
assign g7614 = ((~II12190));
assign g8849 = ((~g8745));
assign g3047 = (g1227&g2306);
assign g1987 = ((~g762));
assign II11342 = ((~g6686));
assign g7277 = (g6772&g731);
assign g8610 = ((~g8483));
assign g2997 = ((~g2135));
assign II15604 = ((~g10148));
assign II17297 = ((~g11369))|((~II17295));
assign gbuf12 = (g1360);
assign g7037 = ((~II11198));
assign g5110 = (g1806&g4618);
assign g3395 = ((~II6601));
assign II13409 = ((~g8141));
assign g6825 = ((~II10873));
assign g7226 = ((~II11464));
assign g10013 = (II15214)|(II15215);
assign g9076 = ((~g8892));
assign II9514 = ((~g5094));
assign II4777 = ((~g18));
assign g10324 = ((~g9317)&(~g10244));
assign g2434 = ((~g1362));
assign II7453 = ((~g3708));
assign g6788 = (g287&g5876);
assign g2237 = ((~g713));
assign II14888 = ((~g9454));
assign g5838 = (g5612)|(g4866);
assign g7887 = ((~g7693));
assign g3423 = (II6630&II6631);
assign II7173 = ((~g2644));
assign II9129 = ((~g4892));
assign II8591 = ((~g501))|((~II8589));
assign g6522 = (g5744)|(g4994);
assign g9391 = ((~g9010)&(~g9240)&(~g9223)&(~II14602));
assign g11184 = ((~II16953));
assign g3371 = ((~g2837));
assign g9679 = ((~g9452));
assign g5593 = ((~II9013));
assign g8872 = ((~II14188));
assign II16735 = ((~g10855));
assign g11396 = ((~II17231));
assign g4904 = (g1850&g4243);
assign II14612 = ((~g9204))|((~g611));
assign II12002 = ((~g7082))|((~g153));
assign g6305 = ((~II10174));
assign II16072 = ((~g845))|((~g10373));
assign g4051 = ((~II7166));
assign II16492 = ((~g10773));
assign g5173 = (g3094&g4676);
assign g3980 = ((~g3121));
assign g4104 = ((~g3215))|((~g3247))|((~g2439))|((~g3200));
assign g5736 = ((~II9296));
assign g9556 = ((~II14701));
assign II17692 = ((~g11596));
assign g10391 = ((~g10313));
assign g6869 = ((~II10949));
assign II12505 = ((~g7728));
assign g7728 = ((~II12369));
assign g8889 = (g8844)|(g8756);
assign g10351 = ((~II15817));
assign g8869 = ((~II14179));
assign g9607 = (g12&g9274);
assign II8605 = ((~g4259))|((~II8604));
assign g4202 = ((~II7423));
assign g6516 = (g5993&g3097);
assign g11405 = ((~II17258));
assign g8009 = ((~II12849));
assign g10064 = ((~II15290));
assign II13636 = ((~g8357));
assign g7721 = (g736&g7237);
assign g8235 = ((~g7967));
assign g9892 = ((~II15079));
assign II13043 = ((~g8055));
assign g4464 = ((~II7829));
assign g4907 = ((~II8278));
assign II17450 = ((~g11450));
assign II6288 = ((~g2091))|((~II6287));
assign g4229 = (g999&g3914);
assign g5858 = ((~II9475));
assign g3008 = ((~g2444))|((~g878));
assign II6110 = ((~g2205))|((~II6109));
assign II14279 = ((~g1828))|((~II14277));
assign g2261 = ((~g1713));
assign II14540 = ((~g9310));
assign II11008 = ((~g6795));
assign g11490 = ((~II17486))|((~II17487));
assign g6424 = ((~g6140));
assign g2610 = ((~II5731));
assign g6221 = (g782&g5598);
assign g6680 = ((~II10643));
assign II16252 = ((~g10515));
assign g6386 = ((~II10282));
assign g7672 = ((~II12293));
assign g10629 = ((~g10583));
assign g9857 = (g9734&g9569);
assign II13102 = ((~g7928));
assign g4994 = (g1504&g4640);
assign g5644 = ((~II9093));
assign g8724 = (g8606&g7910);
assign g5264 = (g1095&g4763);
assign g9352 = ((~II14561));
assign II7345 = ((~g4050));
assign g8344 = ((~II13412));
assign g6242 = ((~II9995));
assign g5122 = ((~g4682));
assign II16273 = ((~g10559));
assign g11056 = ((~g10950));
assign g10423 = ((~g10290)&(~g4620));
assign II8340 = ((~g4804));
assign II5960 = ((~g2239));
assign II9669 = ((~g5426));
assign II11921 = ((~g6904));
assign II6989 = ((~g2760))|((~II6988));
assign g6068 = (g5220)|(g4497);
assign g5503 = ((~g4515));
assign g6449 = ((~g6172));
assign II4961 = ((~g254));
assign II5264 = ((~g456))|((~II5263));
assign g5762 = (g5178)|(g5186);
assign g9590 = (g895&g8995);
assign g9896 = (g9883&g9624);
assign g8156 = ((~II13051));
assign g6440 = ((~g6150));
assign II5821 = ((~g2101));
assign g10800 = (g6245)|(g10772);
assign II13250 = ((~g8148))|((~II13248));
assign g5678 = ((~II9191));
assign g2233 = ((~II5224));
assign g10553 = ((~II16220));
assign II10388 = ((~g5830));
assign g6933 = ((~II11061));
assign II6851 = ((~g2937));
assign g7270 = ((~II11515));
assign g8824 = ((~g8502))|((~g8501))|((~g8739));
assign g7341 = ((~II11671));
assign II10195 = ((~g6116));
assign g7203 = (g6640)|(g6058);
assign II12009 = ((~g6915));
assign g4254 = ((~g4013));
assign g10584 = ((~g10522));
assign II7817 = ((~g3399));
assign g2793 = ((~g2276));
assign II12529 = ((~g7589));
assign II7315 = ((~g2891));
assign II7829 = ((~g3425));
assign g6187 = (g5569&g2340);
assign II15196 = ((~g9974));
assign g7718 = (g709&g7221);
assign g9965 = (g9955&g9536);
assign II7847 = ((~g3435));
assign II11626 = ((~g7042));
assign II15635 = ((~g10185));
assign g5661 = ((~II9144));
assign g8607 = (g8406)|(g8554);
assign g9958 = ((~II15157));
assign g11158 = (g309&g10935);
assign II7625 = ((~g4164));
assign g6574 = ((~II10514));
assign g5801 = ((~g5320));
assign II12971 = ((~g8039));
assign II16080 = ((~g849))|((~II16079));
assign g4299 = ((~g4144));
assign g8952 = ((~II14309));
assign II14918 = ((~g9535));
assign II9737 = ((~g5258));
assign II14306 = ((~g8812));
assign II11728 = ((~g7010));
assign g8475 = ((~g8314));
assign g10634 = (g10604&g3829);
assign II12075 = ((~g7098))|((~II12074));
assign II16175 = ((~g10488));
assign II12133 = ((~g6870));
assign II13901 = ((~g8520))|((~II13900));
assign g6040 = ((~II9655));
assign II6754 = ((~g2906));
assign II14136 = ((~g8775));
assign g6311 = ((~II10192));
assign II12751 = ((~g7626));
assign II5271 = ((~g70));
assign g11624 = (g11595)|(g11571);
assign g8323 = ((~II13351));
assign g11448 = ((~II17394))|((~II17395));
assign II10305 = ((~g6180));
assign g7403 = ((~II11783));
assign g4322 = ((~II7593));
assign g4877 = (g243&g3946);
assign II6590 = ((~g3186));
assign II12029 = ((~g6922));
assign II15241 = ((~g10013));
assign g2122 = ((~II5044));
assign g7419 = ((~g7206));
assign II10753 = ((~g5814));
assign g4953 = ((~II8324));
assign g5044 = (g4348&g1918);
assign g9106 = ((~II14439));
assign g7376 = ((~II11756));
assign g9850 = (g9726&g9560);
assign II12081 = ((~g6934));
assign g5220 = (g1083&g4729);
assign g8721 = ((~g8582));
assign II16808 = ((~g10906));
assign II10027 = ((~g5751));
assign II9202 = ((~g4915));
assign g5511 = ((~II8934));
assign g11180 = ((~II16941));
assign II5036 = ((~g1019))|((~II5034));
assign g11289 = ((~II17070));
assign g6438 = (g5853&g5797);
assign II14045 = ((~g8603));
assign g7126 = ((~II11367));
assign II16742 = ((~g10857));
assign g8592 = ((~II13837));
assign g8579 = ((~II13822));
assign g7742 = (g7217)|(g6743);
assign g8793 = (g8644&g8723);
assign g8574 = (g5679)|(g7853)|(g8465);
assign g6210 = ((~g5205));
assign g5392 = ((~g3369)&(~g4258));
assign g7324 = ((~II11620));
assign g2511 = (g461&g456);
assign g2499 = (II5570)|(II5571);
assign II17281 = ((~g11360))|((~g11357));
assign g10298 = (g8892&g10214);
assign g2518 = ((~g590));
assign g8438 = ((~II13612));
assign g9804 = ((~II14939));
assign g4719 = ((~g3586));
assign g10479 = ((~II16059))|((~II16060));
assign II17344 = ((~g11369));
assign g7420 = ((~II11804));
assign II11817 = ((~g7246));
assign g6342 = (g293&g5886);
assign g5090 = (g1781&g4592);
assign g11204 = (g971&g11083);
assign g9554 = ((~II14697));
assign g9409 = (g1721&g9052);
assign g8442 = ((~II13624));
assign II10733 = ((~g6099));
assign g2909 = ((~II6080));
assign g11373 = ((~II17198));
assign II6055 = ((~g2569));
assign g11434 = ((~II17353));
assign II9461 = ((~g4940));
assign g7098 = ((~II11333));
assign II15344 = ((~g10025));
assign g6165 = ((~g5446));
assign g6911 = (g6342)|(g5681);
assign II12520 = ((~g7415));
assign g7583 = ((~II12068))|((~II12069));
assign II17112 = ((~g11227));
assign g9616 = ((~g9010)&(~g9240)&(~g9223)&(~II14751));
assign g7210 = ((~II11440));
assign g10809 = (g4811&g10754);
assign g6265 = ((~II10054));
assign g2075 = ((~II4883));
assign II9677 = ((~g5190));
assign II10996 = ((~g6786));
assign g7899 = ((~II12683));
assign g8174 = (g5284&g7853);
assign II12108 = ((~g135))|((~II12106));
assign g8969 = ((~II14340));
assign g2820 = ((~II5926));
assign II7593 = ((~g4142));
assign g5654 = ((~II9123));
assign g6359 = (g281&g5898);
assign II13224 = ((~g8261));
assign g5722 = (g1598&g5144);
assign g7336 = ((~II11656));
assign g4588 = ((~g3440))|((~g2745));
assign II11797 = ((~g6852));
assign II14989 = ((~g9813));
assign II6762 = ((~g1448))|((~II6760));
assign g9781 = ((~g9392)&(~g9367));
assign II7357 = ((~g4077));
assign II8308 = ((~g4443));
assign II12339 = ((~g7054));
assign g7218 = (g6655)|(g6070);
assign g10191 = ((~II15551));
assign g7348 = ((~II11692));
assign g10711 = (g5547)|(g10690);
assign g8785 = ((~II14090));
assign II6102 = ((~g2240));
assign II16787 = ((~g10896));
assign II16805 = ((~g10904));
assign II10159 = ((~g5936));
assign g5878 = ((~g5309));
assign g11352 = ((~II17173));
assign II7996 = ((~g3462));
assign II13586 = ((~g8356));
assign II12538 = ((~g7658));
assign g3981 = ((~II7118));
assign g10903 = ((~g10809));
assign g11255 = (g456&g11075);
assign II14958 = ((~g9767));
assign II9305 = ((~g4970));
assign g8775 = (g8628&g5151);
assign g3284 = (g2531&g677);
assign g3330 = ((~II6507));
assign g8604 = ((~g8479));
assign g6625 = (g1218&g6178);
assign g8713 = ((~g8684));
assign II17493 = ((~g11475))|((~II17492));
assign g10302 = ((~II15717))|((~II15718));
assign g8760 = ((~g8670));
assign g3266 = ((~II6436));
assign II10060 = ((~g5752));
assign II16373 = ((~g10593));
assign II7793 = ((~g3783));
assign g5759 = ((~II9341));
assign g2108 = ((~II4992));
assign g5740 = ((~II9302));
assign g11606 = (g11585)|(g11556);
assign g2843 = ((~II5963));
assign g6954 = ((~II11100));
assign g6840 = (g248&g6596);
assign g8110 = ((~g7996));
assign g8417 = (g8246)|(g7721);
assign g6862 = ((~g6720));
assign II8752 = ((~g1125))|((~II8750));
assign g11189 = (g5616&g11064);
assign g6566 = ((~g5791));
assign g4183 = ((~II7366));
assign g8688 = ((~g8507));
assign g2399 = ((~g605));
assign g9882 = ((~g9742)&(~g9536)&(~g9563)&(~II15057));
assign II15814 = ((~g10202));
assign g5095 = ((~II8465));
assign g8306 = ((~II13290));
assign II17773 = ((~g11650));
assign g9712 = (g1528&g9490);
assign g7901 = ((~g7712));
assign g4346 = ((~II7625));
assign g2902 = ((~II6061));
assign g2226 = ((~g86));
assign g10291 = ((~g10247)&(~g3113));
assign g2958 = ((~II6163));
assign II15036 = ((~g9721));
assign g11588 = (g1330&g11547);
assign II13400 = ((~g8236));
assign g4834 = (g219&g3946);
assign g8407 = ((~II13522))|((~II13523));
assign II6777 = ((~g2892))|((~g650));
assign g3906 = ((~g3015));
assign II11770 = ((~g7202));
assign g11201 = (g11152)|(g11011);
assign II10979 = ((~g6565));
assign g2364 = ((~g611));
assign II15353 = ((~g10007));
assign g10821 = ((~II16531));
assign g11210 = (g11078&g4515);
assign g11319 = ((~II17116));
assign II7336 = ((~g3997));
assign g2382 = ((~g599));
assign g9772 = ((~g9432));
assign g10288 = ((~II15688));
assign II11593 = ((~g6830));
assign g2390 = ((~II5475));
assign g9704 = (g9385)|(g9605)|(II14835);
assign II15763 = ((~g10244));
assign II17393 = ((~g11415))|((~g11414));
assign g6128 = ((~II9829));
assign g6283 = ((~II10108));
assign II16184 = ((~g10484));
assign g8366 = (g8199&g7265);
assign g3416 = ((~g3144));
assign g8056 = ((~g7671));
assign II12120 = ((~g7106));
assign g3353 = ((~g3121));
assign g4216 = ((~II7465));
assign II17252 = ((~g11343));
assign g2603 = ((~II5710));
assign II15592 = ((~g10163));
assign g6640 = (g5281&g5801);
assign g3530 = ((~II6715))|((~II6716));
assign g3479 = ((~g2655));
assign g10663 = (g10237)|(g10581);
assign g8772 = (g8627&g5151);
assign gbuf7 = (g1955);
assign II10822 = ((~g6584));
assign g6794 = (g5819&g4415);
assign II7369 = ((~g4051));
assign g6052 = ((~g5426));
assign g11590 = (g2274&g11561);
assign g9822 = ((~II14967));
assign g3811 = ((~II7029));
assign II7852 = ((~g3438));
assign g5697 = ((~II9232));
assign g11149 = (g324&g10930);
assign g7060 = (g6739&g5521);
assign g11392 = (g11278&g7914);
assign g9763 = ((~II14906));
assign g10928 = ((~g10827));
assign g8957 = (g8081&g6368&g8828);
assign g4525 = ((~g3880));
assign g2883 = ((~II6037));
assign g10460 = ((~II15971));
assign g4987 = (g1440&g4682);
assign g11277 = (g4920&g11199);
assign g2004 = ((~II4820));
assign II9349 = ((~g5515));
assign g8378 = ((~II13482));
assign g4638 = ((~g3354));
assign II6498 = ((~g2958));
assign g6527 = ((~II10445));
assign g7891 = (g7471&g7028);
assign g11245 = ((~g11112));
assign II11115 = ((~g6462));
assign g8071 = (g691&g7826);
assign g3386 = ((~g3144));
assign g8842 = (g8607&g8707);
assign g10033 = ((~II15235));
assign II5992 = ((~g2195));
assign g7992 = ((~g7011))|((~g7574))|((~g6984))|((~g6974));
assign II7909 = ((~g3387));
assign g7806 = ((~II12583));
assign II13867 = ((~g8523))|((~g1403));
assign g3693 = ((~g2920));
assign II5053 = ((~g1188));
assign g6091 = ((~II9744));
assign II5916 = ((~g2217));
assign g8990 = ((~II14391));
assign g11597 = (g11576&g5446);
assign II9056 = ((~g4753));
assign g4640 = (g3348)|(g3563)|(g1527);
assign g11101 = (g857&g10950);
assign g11037 = ((~II16772));
assign g3362 = ((~II6546));
assign II12547 = ((~g7673));
assign g6205 = (g1515&g5151);
assign II9822 = ((~g5219));
assign g11314 = (g11224)|(g11102);
assign II11279 = ((~g305))|((~II11278));
assign g2454 = ((~II5549));
assign g2459 = ((~g1645)&(~g1642)&(~g1651)&(~g1648));
assign g7621 = (g5108)|(g6994);
assign II14509 = ((~g8926));
assign g9506 = ((~g9052)&(~g9030));
assign g6778 = ((~g5987));
assign II11719 = ((~g7029));
assign g11217 = (g11144)|(g11005);
assign g6289 = ((~II10126));
assign g9908 = (g9890&g9782);
assign g6895 = (g6776)|(g4875);
assign g7813 = ((~II12604));
assign II11467 = ((~g6488));
assign g4232 = ((~II7487));
assign II6686 = ((~g3015));
assign g6583 = ((~II10535));
assign g9931 = (g8931)|(g9900);
assign II11217 = ((~g6529));
assign g6591 = ((~II10553));
assign g6182 = ((~g5446));
assign II10165 = ((~g5948));
assign g11503 = ((~II17528));
assign II8031 = ((~g3540));
assign II12326 = ((~g7246));
assign II13812 = ((~g8519));
assign g7977 = ((~II12779));
assign II5935 = ((~g2174));
assign II8730 = ((~g1117))|((~II8728));
assign II7295 = ((~g3260));
assign II7006 = ((~g2912));
assign II6480 = ((~g2462));
assign g7195 = ((~II11417));
assign g9664 = (g1191&g9125);
assign g3775 = ((~II7002));
assign g8317 = ((~II13335));
assign II14182 = ((~g8788));
assign g5980 = ((~II9594));
assign g8040 = (g7523&g5128);
assign II13109 = ((~g7981));
assign g10346 = ((~II15804));
assign II5203 = ((~g369))|((~II5202));
assign II8039 = ((~g3506));
assign g7356 = ((~II11716));
assign g11328 = (g11299)|(g11168);
assign g9692 = (g272&g9432);
assign II7378 = ((~g4067));
assign g3763 = ((~II6968));
assign g2303 = ((~II5342))|((~II5343));
assign g7608 = ((~II12174));
assign g7041 = ((~g6427));
assign g7526 = (g7148&g2868);
assign g6059 = (g5211)|(g4489);
assign II13290 = ((~g8254));
assign g9349 = ((~II14552));
assign g10449 = (g10420&g3345);
assign g10205 = ((~g10176));
assign g7932 = ((~g7395))|((~g6847))|((~g7279))|((~g7273));
assign g4362 = ((~II7651));
assign g11078 = ((~II16847));
assign g5659 = ((~II9138));
assign II15302 = ((~g10007));
assign II15479 = ((~g10091));
assign g9732 = ((~II14873));
assign II9371 = ((~g5075));
assign g10621 = ((~II16298));
assign II9043 = ((~g4786));
assign g11269 = (g11196)|(g11031);
assign g7987 = ((~g7011))|((~g6995))|((~g7562))|((~g6974));
assign g6763 = (g5802&g4381);
assign g10802 = ((~II16510));
assign g4604 = (g3056&g3753&g2325);
assign g10442 = (g10311&g2135);
assign g8116 = ((~II12971));
assign II7291 = ((~g3212));
assign g10489 = (g4961)|(g10367);
assign g7042 = ((~II11211));
assign II11587 = ((~g6828));
assign g3432 = ((~g3144));
assign g6132 = ((~II9833));
assign g5474 = ((~II8889));
assign g9760 = ((~g9454));
assign II5940 = ((~g2175));
assign g5852 = (g5632)|(g4883);
assign g4008 = (g2689&g2276);
assign g9860 = (g1598&g9775);
assign II11091 = ((~g6657));
assign g5754 = ((~II9332));
assign g9754 = (g9173)|(g9511);
assign g3425 = (g2895)|(g2910);
assign II10135 = ((~g6249));
assign g6397 = ((~II10299));
assign II7716 = ((~g3751));
assign g6689 = ((~g5830));
assign II13203 = ((~g8196));
assign II8418 = ((~g4794));
assign II5867 = ((~g2105))|((~II5865));
assign g7775 = ((~II12490));
assign g11581 = (g1308&g11539);
assign g4377 = ((~II7694));
assign g8094 = ((~g7987));
assign g8076 = ((~II12930));
assign g11510 = ((~II17549));
assign g10555 = (g4103)|(g10504);
assign II16920 = ((~g11084));
assign g6178 = ((~g4977));
assign II5295 = ((~g794))|((~g798));
assign g8389 = (g6091&g8225);
assign g5212 = (g1255&g4726);
assign g4193 = ((~II7396));
assign II12904 = ((~g7985));
assign g9887 = ((~II15068));
assign g10589 = ((~II16252));
assign g5690 = (g1567&g5112);
assign II5613 = ((~g1284))|((~II5611));
assign g7309 = ((~II11575));
assign II13197 = ((~g8186));
assign II14961 = ((~g9769));
assign II14779 = (g8995)|(g9205)|(g9192);
assign II7240 = ((~g2824));
assign g3537 = ((~g3164));
assign II9875 = ((~g5278));
assign g10368 = ((~g10342)&(~g3463));
assign II13266 = ((~g1909))|((~II13265));
assign II5025 = ((~g1275))|((~II5023));
assign g7737 = ((~II12388));
assign g5034 = ((~g3524)&(~g4593));
assign g2339 = ((~II5399));
assign II5672 = ((~g569));
assign g10283 = ((~g10166));
assign g4498 = (g1145&g3940);
assign g7637 = ((~II12251));
assign g3996 = ((~g3144));
assign g11348 = ((~g11276));
assign g3519 = ((~g3164));
assign II9023 = ((~g4727));
assign g7706 = ((~II12335));
assign g2652 = ((~g2008));
assign g11042 = ((~II16787));
assign g11384 = ((~II17209));
assign g2069 = ((~II4869));
assign g10500 = (g4157)|(g10442);
assign g7730 = (g7260&g2347);
assign g11175 = (g501&g11112);
assign g4879 = ((~g3292)&(~g2593)&(~g3784)&(~g2579));
assign g6154 = ((~II9875));
assign g4794 = ((~II8164));
assign g8615 = (g8413)|(g8557);
assign II10144 = ((~g5689));
assign g2255 = ((~II5276));
assign II7559 = ((~g4116));
assign g6081 = ((~g4977));
assign II15807 = ((~g10284));
assign g4191 = ((~II7390));
assign g7046 = (g5892&g6570);
assign g11555 = (g2695&g11519);
assign g10161 = ((~II15479));
assign II17331 = ((~g11357));
assign II9365 = ((~g5392));
assign II15565 = ((~g10101));
assign II9539 = ((~g5354));
assign II8535 = ((~g4340));
assign II5342 = ((~g315))|((~II5341));
assign g5866 = ((~g5361));
assign II13877 = ((~g8535))|((~II13876));
assign II13051 = ((~g8060));
assign II13436 = ((~g8187));
assign g7473 = ((~g7148));
assign II17108 = ((~g11225));
assign II15057 = (g7853)|(g9680)|(g9624)|(g9785);
assign g8674 = ((~II13959));
assign g8701 = (g7597&g8582);
assign g10156 = ((~II15464));
assign g2216 = ((~g41));
assign g6348 = (g296&g5891);
assign g6203 = ((~g5446));
assign II10659 = ((~g6038));
assign g6482 = ((~II10412));
assign II17616 = ((~g11561));
assign g5598 = (g778&g4824);
assign g9746 = ((~g9454)&(~g9274)&(~g9292));
assign g98 = ((~II4783));
assign g8177 = ((~II13077))|((~II13078));
assign g8748 = (g7670&g8656);
assign II7639 = ((~g3722));
assign g8656 = ((~II13941));
assign II14252 = ((~g8783));
assign g5591 = (g1615&g4514);
assign g10354 = ((~II15826));
assign g5700 = ((~II9237));
assign II15994 = ((~g2677))|((~II15992));
assign II8282 = ((~g4770));
assign g11084 = ((~II16863));
assign g4262 = ((~g4013));
assign g8754 = (g7420&g8667);
assign II15082 = ((~g9719));
assign II16601 = ((~g10806));
assign g3098 = (g2331&g2198);
assign g6442 = ((~II10362));
assign II14112 = ((~g8777));
assign II5922 = ((~g2170));
assign g8420 = ((~II13574));
assign II12436 = ((~g7659));
assign g9653 = (g1185&g9125);
assign g5830 = ((~II9446));
assign g10643 = (g10624)|(g7736);
assign g7466 = (g7148&g2821);
assign g2007 = ((~g936));
assign II8662 = ((~g4286))|((~g476));
assign g5081 = ((~II8449));
assign II10963 = ((~g6793));
assign II5591 = ((~g1696))|((~g1703));
assign g5032 = ((~II8403));
assign g6463 = (g5052&g6210);
assign g6880 = (g4816&g6562);
assign g11085 = (g312&g10897);
assign g2807 = ((~g22)&(~g2320));
assign II16956 = ((~g11096));
assign g6088 = (g5260)|(g4522);
assign II17503 = ((~g11475))|((~g7603));
assign g4504 = ((~II7899));
assign g8194 = (g5168)|(g7940);
assign g9939 = (g9918&g9367);
assign g5671 = ((~II9174));
assign g10065 = ((~II15293));
assign g8627 = ((~II13887))|((~II13888));
assign II16160 = (g10394)|(g10392)|(g10482)|(g10481);
assign g7687 = ((~II12318));
assign g8963 = (g8056&g6368&g8849);
assign g10111 = ((~II15347));
assign g5481 = ((~II8900));
assign II10183 = ((~g6108));
assign g2861 = ((~II6001));
assign g3086 = ((~g2276));
assign g2021 = ((~g1341));
assign II9544 = ((~g5024));
assign g2028 = ((~g1703));
assign g11076 = ((~II16843));
assign g8929 = (g8095&g6368&g8828);
assign II6952 = ((~g2867));
assign g10458 = ((~II15965));
assign g7627 = ((~II12223));
assign II15332 = ((~g10001));
assign g10327 = ((~II15771));
assign g6073 = ((~II9712));
assign g10534 = ((~II16169));
assign g3337 = ((~g2745));
assign II11836 = ((~g7220));
assign g8922 = (g8822)|(g8736);
assign g7384 = (g7088)|(g6618);
assign II15716 = ((~g10231))|((~g10229));
assign g3707 = ((~g2920));
assign g6750 = ((~II10759));
assign g11423 = ((~II17324));
assign g6647 = (g5288&g5808);
assign g10775 = ((~II16461));
assign g7183 = (g6623)|(g6046);
assign g5072 = ((~II8442));
assign g3877 = ((~II7064));
assign g10041 = ((~II15250));
assign g11408 = ((~II17265));
assign II7435 = ((~g3459));
assign g5169 = ((~g4596));
assign g6694 = ((~II10663));
assign g4286 = ((~g3800)&(~g2593)&(~g3784)&(~g2579));
assign g2946 = ((~II6133));
assign g6576 = (g5762&g5503);
assign g5039 = ((~II8418));
assign g7782 = ((~II12511));
assign g11112 = ((~II16897));
assign g2629 = ((~g2001));
assign g7029 = ((~II11180));
assign g2205 = ((~II5165))|((~II5166));
assign g7773 = ((~II12484));
assign g3814 = ((~g3228));
assign g9852 = (g9728&g9563);
assign g9943 = (g9923&g9367);
assign II16017 = ((~g2695))|((~II16015));
assign g8291 = ((~II13227));
assign g5887 = ((~II9510));
assign g1964 = ((~g114));
assign II16065 = ((~g10428))|((~g2765));
assign g7335 = ((~II11653));
assign g9430 = (g1759&g9030);
assign g8569 = ((~II13800));
assign g11264 = (g11188)|(g11026);
assign g9697 = (g9665)|(g9606)|(II14822);
assign II9276 = ((~g5241));
assign g7231 = (g6673)|(g6087);
assign g4079 = (g2765&g2276);
assign g3521 = ((~g3164));
assign II12427 = ((~g7636));
assign g6039 = ((~II9652));
assign g11638 = ((~II17724));
assign II8611 = ((~g4562));
assign II4886 = ((~g257));
assign g10529 = (II16160)|(II16161);
assign II14973 = ((~g9733));
assign g10612 = ((~II16286));
assign g4440 = ((~g4130));
assign g8330 = ((~II13370));
assign g9418 = (g1741&g9052);
assign g10798 = (g6217)|(g10768);
assign g4872 = ((~II8211));
assign g6801 = ((~II10813));
assign g5285 = ((~g4355));
assign II4986 = ((~g999))|((~II4985));
assign g11098 = (g849&g10950);
assign g9802 = ((~g9490));
assign g3752 = ((~II6947));
assign g2914 = ((~II6091));
assign g2986 = ((~II6220));
assign g3528 = ((~g3164));
assign g5817 = ((~II9427));
assign II9016 = ((~g4722));
assign g10856 = (g6083)|(g10737);
assign g4971 = (g1419&g4682);
assign g5532 = (g1681&g4307);
assign II16236 = ((~g10535));
assign g9365 = (g1321&g9151);
assign g8339 = ((~II13397));
assign II10231 = ((~g6111));
assign g4771 = (g496&g3416);
assign g4801 = (g516&g3439);
assign II5248 = ((~g1110));
assign II7803 = ((~g3820));
assign II11915 = ((~g6935))|((~II11914));
assign g6251 = ((~II10012));
assign g9270 = ((~II14485));
assign g3941 = ((~g3015));
assign II5430 = ((~g916));
assign II6037 = ((~g2560));
assign g5225 = ((~II8663))|((~II8664));
assign g3113 = ((~II6343));
assign II6815 = ((~g2755));
assign g5796 = (g1564&g5252);
assign II8750 = ((~g4613))|((~g1125));
assign g2530 = ((~II5641));
assign g2731 = ((~II5789));
assign II7478 = ((~g3566));
assign g2259 = ((~II5292));
assign g6732 = ((~II10729));
assign g7954 = (g2874&g7512);
assign II6022 = ((~g2258));
assign g8818 = (g7955)|(g8733);
assign II12106 = ((~g7113))|((~g135));
assign II5283 = ((~g758))|((~II5282));
assign g3943 = ((~g2779));
assign g3736 = ((~II6924));
assign g6843 = ((~II10901));
assign g8358 = ((~II13454));
assign II14216 = ((~g8826))|((~g605));
assign g3688 = (g3144)|(g2454);
assign II14684 = ((~g9124));
assign g8203 = (g7453)|(g7999);
assign II6186 = ((~g2511))|((~g466));
assign g11610 = (g11589)|(g11560);
assign g10277 = ((~II15675));
assign g4082 = ((~II7213));
assign g2347 = ((~g1945));
assign II11937 = ((~g1458))|((~II11935));
assign g9173 = (g8968&g6674);
assign g7541 = (g7075&g3109);
assign g9721 = (g9413&g4785);
assign II14903 = ((~g9507));
assign g7548 = ((~II11981))|((~II11982));
assign g4765 = (g491&g3405);
assign g5508 = ((~II8929));
assign g4425 = ((~II7771));
assign II4942 = ((~g396))|((~II4941));
assign II14203 = ((~g8825))|((~II14202));
assign II15545 = ((~g10075));
assign g9340 = ((~II14525));
assign II15263 = ((~g9995));
assign g3698 = (g3121)|(g2480);
assign II15968 = ((~g10408));
assign II15878 = ((~g10359))|((~g2719));
assign g5826 = ((~II9440));
assign g3247 = ((~g1828))|((~g2564))|((~g2571));
assign g9844 = (g9714&g9522);
assign g3582 = ((~g3164));
assign g8858 = ((~g8743));
assign g11179 = ((~II16938));
assign II16859 = ((~g10911));
assign g9819 = ((~II14958));
assign II10643 = ((~g6026));
assign g2168 = ((~II5111));
assign II16553 = ((~g10754));
assign g8484 = ((~g8336));
assign II6968 = ((~g2881));
assign II15253 = ((~g9987));
assign g6323 = (g1235&g5949);
assign II14424 = ((~g8945));
assign g10431 = ((~g10328));
assign g2745 = ((~II5809));
assign g8935 = (g8106&g6778&g8849);
assign II7280 = ((~g3208));
assign II17146 = ((~g11305));
assign g4530 = ((~II7935));
assign g7824 = (g1932&g7479);
assign g3635 = ((~II6812));
assign g10541 = ((~II16190));
assign g9974 = (II15176)|(II15177);
assign II17387 = ((~g11438));
assign g6134 = ((~II9839));
assign II5710 = ((~g2431));
assign II13531 = ((~g8253))|((~II13529));
assign II7061 = ((~g3050));
assign g10168 = ((~II15500));
assign II14040 = ((~g8649));
assign g11292 = (g11252&g4250);
assign g5249 = (g1089&g4747);
assign g7561 = ((~II12015));
assign g10426 = ((~g10294)&(~g4620));
assign g2643 = ((~g1989));
assign g9689 = (g263&g9432);
assign g4913 = ((~II8285));
assign g4593 = ((~II8004));
assign g5479 = (g1845&g4243);
assign g5732 = (g1604&g5176);
assign g8429 = (g8385)|(g8069);
assign g4351 = ((~II7630));
assign g4520 = ((~II7923));
assign g5402 = ((~II8842));
assign g4256 = ((~g3664));
assign g4163 = ((~II7308));
assign g7302 = (g7141)|(g6328);
assign g7007 = ((~II11146));
assign g8512 = ((~g3723))|((~g8366));
assign g8519 = ((~II13726));
assign g4935 = ((~g4420));
assign II11207 = ((~g6524));
assign g2772 = ((~g2508));
assign g6275 = ((~II10084));
assign II9102 = ((~g5586));
assign g11412 = ((~II17277));
assign g11505 = ((~II17534));
assign g11592 = (g3717&g11561);
assign II8827 = ((~g4477));
assign II13248 = ((~g1891))|((~g8148));
assign g2617 = ((~g1997));
assign g4315 = ((~g3863));
assign g9816 = ((~g9490));
assign g3744 = ((~g3307));
assign II5357 = (g1265)|(g1260)|(g1255)|(g1250);
assign II6310 = (g2396&g2407&g2421&g2435);
assign g7242 = (g6693)|(g6098);
assign g10088 = ((~II15317));
assign g2363 = ((~II5441));
assign II16427 = (g10683)|(g10608)|(g10604);
assign g8387 = (g6086&g8220);
assign g6106 = ((~II9773));
assign g4734 = ((~g3586));
assign g5842 = (g5618)|(g4870);
assign g6326 = (g1250&g5949);
assign g5663 = ((~II9150));
assign g2047 = ((~g1857));
assign g8128 = ((~II12993));
assign g8002 = ((~II12832));
assign g3038 = ((~g1982));
assign g10875 = ((~II16595));
assign II11908 = ((~g6967))|((~II11907));
assign g4251 = ((~g3292)&(~g3793)&(~g3784)&(~g2579));
assign II9147 = ((~g5011));
assign g7260 = (g6752&g2345);
assign II9194 = ((~g5236));
assign II5892 = ((~g750))|((~II5891));
assign II6767 = ((~g2914));
assign g6272 = ((~II10075));
assign II12114 = ((~g7093))|((~II12113));
assign g10736 = (g10658&g4840);
assign g8264 = (g7879)|(g3389);
assign g4780 = ((~g3440));
assign II5005 = ((~g421))|((~g312));
assign g4727 = (g386&g3364);
assign II15736 = ((~g10258));
assign g3977 = ((~II7112));
assign g4487 = (g1718&g3911);
assign II17246 = ((~g11341));
assign II11665 = ((~g7038));
assign II14415 = ((~g8940));
assign g8015 = ((~II12857));
assign II6040 = ((~g2216));
assign g6727 = ((~g5997));
assign g10691 = ((~II16360));
assign II5865 = ((~g2107))|((~g2105));
assign II15443 = ((~g10122))|((~II15441));
assign II15607 = ((~g10149))|((~g10144));
assign g9840 = (g9704&g9747);
assign g8433 = (g8399)|(g8073);
assign g2325 = ((~g611))|((~g617));
assign g4275 = ((~g3664));
assign II13969 = ((~g8451));
assign g7063 = (g5903&g6582);
assign II4928 = ((~g391))|((~g321));
assign II10549 = ((~g6184));
assign g10898 = (g4220)|(g10777);
assign g10973 = ((~II16720));
assign g8283 = (g8098)|(g7820);
assign g8949 = (g8255&g6368&g8828);
assign II15775 = ((~g10253));
assign g7437 = ((~II11829));
assign II13415 = ((~g8144));
assign g11321 = (g11230)|(g11105);
assign II11155 = ((~g6470));
assign g5415 = ((~II8848));
assign II6007 = ((~g2199));
assign g10706 = (g10567&g4840);
assign II16032 = ((~g10368))|((~II16030));
assign II6821 = ((~g3015));
assign g6433 = ((~II10349));
assign g6559 = ((~g5758));
assign g5271 = (g727&g4772);
assign g9724 = (g9409)|(g9419)|(g9615);
assign g10885 = ((~g10809));
assign g3102 = ((~g2482));
assign g9641 = (g913&g9205);
assign g10208 = ((~II15580));
assign II16416 = ((~g10664));
assign II7308 = ((~g3070));
assign g5115 = (g1394&g4572);
assign g7800 = ((~II12565));
assign g5771 = (g1534&g5213);
assign II7384 = ((~g4082));
assign g11308 = (g11218)|(g11098);
assign g7496 = (g7148&g2840);
assign II16467 = ((~g10716))|((~g10518));
assign g2097 = ((~II4935));
assign II9658 = ((~g5150));
assign g8483 = ((~g8332));
assign II9588 = ((~g5114));
assign g4159 = ((~II7300));
assign g3747 = ((~g3015));
assign g6266 = ((~II10057));
assign II10186 = ((~g6110));
assign g8183 = ((~II13102));
assign II13529 = ((~g704))|((~g8253));
assign II5202 = ((~g369))|((~g374));
assign g10242 = ((~II15632));
assign g11211 = (g11058&g5534);
assign II12245 = ((~g7093));
assign II5606 = ((~g1153))|((~II5604));
assign g3544 = ((~g3164));
assign g8589 = ((~II13834));
assign II5126 = ((~g1386))|((~g1389));
assign g10633 = (g10600&g3829);
assign g8450 = ((~II13648));
assign II9132 = ((~g4893));
assign g10098 = ((~II15332));
assign g3880 = (g3186&g2023);
assign II15554 = ((~g10088));
assign g10491 = ((~II16108));
assign g10314 = ((~II15744));
assign g4400 = (g4088&g3829);
assign II11119 = ((~g6461));
assign II13364 = ((~g8221));
assign g4921 = (g2779&g4431);
assign II12999 = ((~g7844));
assign g2635 = ((~g2003));
assign g4475 = ((~II7852));
assign II7390 = ((~g4087));
assign II10081 = ((~g5735));
assign g7764 = ((~II12457));
assign II12235 = ((~g7082));
assign g2276 = (g1765&g1610);
assign II15615 = ((~g10043))|((~g10153));
assign g5586 = ((~II8996));
assign g2170 = ((~g30));
assign g5918 = (g2965&g5292&g4609);
assign g7807 = ((~II12586));
assign g9812 = ((~g9490));
assign g11027 = (g391&g10974);
assign g4230 = (g1095&g3638);
assign g8513 = ((~II13708));
assign g2895 = (g2411&g1678);
assign g2195 = ((~g83));
assign g11542 = ((~g11519));
assign II15290 = ((~g9984));
assign II5098 = ((~g38));
assign g8561 = ((~II13776));
assign II15232 = ((~g9974));
assign g3722 = ((~II6894));
assign g8693 = (g3738&g8509);
assign g10744 = (g10600)|(g10668)|(II16427);
assign g9313 = (g8876&g5708);
assign g7444 = (g7277&g5827);
assign II10729 = ((~g5935));
assign II16439 = ((~g10702));
assign II7264 = ((~g3252));
assign g4894 = ((~II8247));
assign g8551 = ((~g3967))|((~g8390));
assign II5549 = ((~g868));
assign II6904 = ((~g2820));
assign g7240 = (g6687)|(g6095);
assign II11169 = ((~g6481));
assign g4060 = ((~g3144));
assign g9308 = ((~II14499));
assign g10664 = (g10240)|(g10582);
assign g11280 = (g11254)|(g11153);
assign g5291 = ((~g4384));
assign g7958 = (g736&g7697);
assign g11153 = (g3771&g10913);
assign g5810 = (g5588)|(g4823);
assign g11151 = (g327&g10931);
assign II9948 = ((~g1796))|((~II9946));
assign g9865 = (g1607&g9780);
assign g3791 = ((~II7014));
assign g5278 = ((~II8739))|((~II8740));
assign g9662 = (g2094&g9292);
assign g1972 = ((~g461));
assign g7585 = ((~II12081));
assign g8298 = ((~II13249))|((~II13250));
assign g11104 = (g2963&g10937);
assign g9994 = ((~II15196));
assign g5002 = (g1494&g4640);
assign g3214 = ((~II6391));
assign II8716 = ((~g4601))|((~II8715));
assign g3563 = (g3275&g2126);
assign g9735 = (g9649)|(g9651)|(g9384)|(g9361);
assign g6121 = ((~II9816));
assign II5332 = ((~g756));
assign II11638 = ((~g6948));
assign g10235 = ((~g10189));
assign g7501 = ((~II11879));
assign g6823 = (g1368&g6596);
assign II5035 = ((~g1015))|((~II5034));
assign g9614 = (g1197&g9111);
assign II13895 = ((~g1436))|((~II13893));
assign g8880 = ((~II14203))|((~II14204));
assign II8275 = ((~g4351));
assign II13767 = ((~g8417))|((~II13765));
assign g10671 = (g10578&g9431);
assign g4122 = ((~g3291)&(~g2410)&(~g2538));
assign g9587 = (g892&g8995);
assign II8943 = ((~g4585));
assign II17395 = ((~g11414))|((~II17393));
assign g5146 = ((~g4596));
assign II9427 = ((~g4963));
assign g7286 = ((~II11534));
assign g6545 = (g5795)|(g5025);
assign g6903 = ((~II11005));
assign II9886 = ((~g5286));
assign II7194 = ((~g2629));
assign II5198 = ((~g143));
assign g2235 = ((~g96));
assign g2919 = ((~II6102));
assign II8589 = ((~g4251))|((~g501));
assign II8967 = ((~g4482));
assign g11236 = (g5469&g11108);
assign g7630 = ((~II12232));
assign g7876 = (g7609&g3790);
assign g4175 = ((~II7342));
assign g11602 = (g11581)|(g11552);
assign g4962 = (g1651&g4461);
assign II13726 = ((~g8375));
assign II16044 = ((~g833))|((~g10370));
assign g5876 = ((~g5361));
assign g10434 = ((~g10352)&(~g3566));
assign g2011 = ((~g976));
assign g7872 = ((~II12655));
assign g6740 = ((~g6131))|((~g2550));
assign II13086 = ((~g7924));
assign g9516 = (g9151)|(g9125);
assign g9026 = ((~II14415));
assign II15801 = ((~g10282));
assign g5614 = ((~II9040));
assign II13505 = ((~g677))|((~II13504));
assign II8385 = ((~g4238));
assign g3307 = ((~II6480));
assign g2868 = ((~II6010));
assign g9968 = (II15171)|(II15172);
assign g6338 = ((~II10237));
assign g6714 = ((~g5867));
assign g11479 = ((~II17470));
assign g11444 = ((~II17381));
assign g5611 = (g1047&g4382);
assign g9918 = (g9858)|(g9698);
assign II5484 = ((~g1250))|((~g1011));
assign II11578 = ((~g6824));
assign g7294 = (g7068)|(g6320);
assign g5893 = ((~g5106));
assign g2310 = ((~g591))|((~g605));
assign II16843 = ((~g10898));
assign g4870 = (g237&g3946);
assign II7076 = ((~g2985));
assign II16623 = ((~g10858));
assign g7649 = ((~II12258));
assign g2570 = ((~g207));
assign g6759 = (g148&g5919);
assign g6297 = ((~II10150));
assign II8669 = ((~g4831))|((~g814));
assign g8707 = ((~g8671));
assign g4672 = ((~g3501)&(~g2669)&(~g2662)&(~g3479));
assign g8879 = (g8110&g6764&g8858);
assign II15177 = (g9844)|(g9960)|(g9863)|(g9876);
assign g4828 = (g4106&g695);
assign II17377 = ((~g11412));
assign g8101 = (g6208&g7877);
assign g4888 = ((~II8237));
assign II15752 = ((~g10264));
assign II17736 = ((~g11640));
assign II12162 = ((~g7146));
assign II14442 = ((~g8970))|((~g1834));
assign g8328 = ((~II13364));
assign g2249 = ((~g127));
assign II15823 = ((~g10201));
assign g9912 = (g9847)|(g9690);
assign g8813 = (g7943)|(g8726);
assign II5494 = ((~g1690));
assign g8266 = (g7885)|(g3412);
assign II6088 = ((~g2235));
assign g11036 = ((~II16769));
assign II12616 = ((~g7534));
assign g6413 = ((~II10325));
assign II12799 = ((~g7556));
assign II15063 = ((~g9699));
assign II10495 = ((~g6144));
assign g11578 = ((~II17616));
assign g5631 = (g1056&g4416);
assign II6121 = ((~g2121));
assign II16023 = ((~g10426))|((~g2701));
assign II4955 = ((~g401))|((~II4954));
assign II8647 = ((~g4219));
assign II13949 = ((~g8451));
assign g8148 = (g7884)|(g6872);
assign II14090 = ((~g8771));
assign g10563 = ((~g10539)&(~g10322));
assign g2537 = ((~II5646));
assign II12255 = ((~g7203));
assign II10036 = ((~g5701));
assign II15977 = ((~g10411));
assign II11082 = ((~g6749));
assign g6723 = ((~II10716));
assign II5716 = ((~g2068));
assign II11982 = ((~g1482))|((~II11980));
assign II13800 = ((~g8500));
assign g10514 = (g10489&g4580);
assign g9898 = (g9887&g9367);
assign II7536 = ((~g4098));
assign g2640 = ((~g1984));
assign II11198 = ((~g6521));
assign g8744 = ((~g8617))|((~g6509))|((~g6971));
assign II13448 = ((~g8150));
assign II8761 = ((~g4616))|((~g1129));
assign g6921 = ((~II11037));
assign g6257 = ((~II10030));
assign g10142 = ((~II15424));
assign g8840 = ((~g8542))|((~g8541))|((~g8760));
assign g4563 = ((~g3946));
assign g4252 = (g1007&g3914);
assign g11489 = ((~II17482));
assign II11932 = ((~g6908));
assign g7967 = ((~II12765));
assign g10421 = ((~g10331));
assign g6806 = ((~II10828));
assign g4483 = (g336&g3586);
assign II12038 = ((~g6990))|((~g1466));
assign g11571 = (g2018&g11561);
assign II8262 = ((~g4636));
assign g10477 = ((~II16045))|((~II16046));
assign II8880 = ((~g4537));
assign g3501 = ((~g3077));
assign g9618 = (g910&g9205);
assign II12690 = ((~g7555));
assign II5641 = ((~g546));
assign g9710 = (g1586&g9474);
assign II17698 = ((~g11616));
assign g9779 = ((~g9392)&(~g9367));
assign II12825 = ((~g7696));
assign g10149 = ((~II15442))|((~II15443));
assign g7611 = ((~II12183));
assign g8181 = ((~II13096));
assign g4591 = ((~g3829));
assign g4534 = (g363&g3586);
assign g4519 = ((~II7920));
assign II11950 = ((~g6906));
assign g7579 = ((~II12053));
assign g2795 = ((~II5892))|((~II5893));
assign g9890 = ((~II15075));
assign g5803 = (g5575)|(g4820);
assign g11156 = (g333&g10934);
assign g8599 = ((~g8546));
assign g7422 = ((~II11810));
assign g10127 = ((~II15383));
assign II9880 = ((~g5405));
assign II5887 = (g2078&g2083&g166&g2095);
assign II5106 = ((~g435))|((~II5104));
assign g10293 = ((~II15701));
assign g4087 = ((~II7220));
assign g3344 = ((~II6528));
assign g8312 = ((~II13320));
assign g4200 = ((~II7417));
assign II4879 = ((~g256));
assign II16717 = ((~g10779));
assign g11607 = (g11586)|(g11557);
assign g2817 = ((~II5919));
assign II14388 = ((~g8924));
assign II5470 = ((~g999))|((~II5468));
assign g8822 = (g8614&g8752);
assign g11394 = ((~II17225));
assign II6888 = ((~g2960));
assign II15551 = ((~g10080));
assign g8308 = ((~II13301))|((~II13302));
assign g4130 = ((~g3044))|((~g2518));
assign II6094 = ((~g2110));
assign g9719 = (g1543&g9490);
assign g6508 = (g5983&g3096);
assign g2424 = ((~g1690));
assign g2654 = ((~g2012));
assign g9600 = (g904&g9205);
assign g8321 = ((~II13347));
assign g5652 = ((~II9117));
assign g4271 = ((~g3971));
assign g6317 = (g1304&g5949);
assign g7749 = ((~II12412));
assign g5657 = ((~II9132));
assign g4806 = (g3215&g3992&g2493);
assign g6907 = (g6792)|(g5675);
assign g9388 = (g9240)|(g9223);
assign g6163 = (g4572&g5354);
assign II13568 = ((~g8343));
assign II11575 = ((~g6823));
assign II8624 = ((~g4267))|((~g511));
assign II10343 = ((~g6003));
assign g3397 = ((~g2896));
assign g2904 = ((~II6065));
assign g8609 = (g8408)|(g8555);
assign g11354 = ((~II17179));
assign II15432 = ((~g10044))|((~II15430));
assign g11432 = ((~II17347));
assign g2352 = ((~II5430));
assign g7845 = ((~II12634));
assign g4974 = ((~g4502)&(~g3714));
assign g4768 = ((~II8126));
assign II12156 = ((~g6878));
assign II5600 = (g496)|(g491)|(g486)|(g481);
assign g10826 = ((~II16540));
assign g8244 = (g7847&g4336);
assign g7921 = ((~g7463));
assign II13609 = ((~g8312));
assign g5426 = ((~II8869));
assign g2905 = ((~II6068));
assign g7032 = (g2965&g6626&g5292);
assign g10551 = ((~II16214));
assign g5769 = (g2112&g4921&g3818);
assign g8146 = ((~g8033));
assign II13975 = ((~g8588));
assign II17444 = ((~g11446));
assign g6666 = (g5301&g5818);
assign g2514 = (II5599)|(II5600);
assign g4319 = ((~g4144));
assign g2071 = ((~II4873));
assign II5976 = ((~g2186));
assign g3096 = ((~g2482));
assign II7272 = ((~g3253));
assign g4452 = ((~g3365));
assign g6734 = ((~II10733));
assign II10147 = ((~g5697));
assign g3304 = ((~II6468))|((~II6469));
assign II14642 = ((~g9088));
assign g6737 = ((~g6016));
assign g5214 = ((~g4640));
assign g2231 = ((~II5218));
assign g7311 = ((~II11581));
assign g6820 = (g1362&g6596);
assign g4375 = ((~g3638));
assign g8572 = ((~II13809));
assign g1963 = ((~g110));
assign g5204 = (g4838&g2126);
assign II13580 = ((~g8338));
assign g7085 = ((~II11318));
assign g8042 = (g7533&g5128);
assign II9326 = ((~g5320));
assign g8472 = ((~II13666));
assign g4297 = ((~II7563))|((~II7564));
assign II10045 = ((~g5727));
assign II6049 = ((~g2219));
assign g9362 = ((~g9010)&(~g9240)&(~g9223)&(~II14585));
assign g10220 = ((~II15592));
assign II17381 = ((~g11436));
assign g6551 = (g5804)|(g5031);
assign g5572 = ((~II8989));
assign II13991 = ((~g622))|((~II13990));
assign g5042 = ((~g4840));
assign g11206 = ((~II16979));
assign g2874 = ((~II6022));
assign II6898 = ((~g2964));
assign g7923 = ((~g7527));
assign II13048 = ((~g8059));
assign g4761 = ((~g3440));
assign II5304 = ((~g79));
assign g9094 = ((~g8892));
assign g4990 = (g1444&g4682);
assign II5655 = ((~g557));
assign g7994 = ((~g7011))|((~g7574))|((~g6984))|((~g7550));
assign II9981 = ((~g5514));
assign g7035 = ((~II11194));
assign g9921 = (g9862)|(g9703);
assign II17209 = ((~g11289));
assign g2187 = ((~g746));
assign II13382 = ((~g8134));
assign II7743 = ((~g3762));
assign g8179 = ((~II13086));
assign II15500 = ((~g10051));
assign g11054 = ((~g10950));
assign II12248 = ((~g7098));
assign g10719 = (g10303)|(g10666);
assign II9585 = ((~g5241));
assign II8854 = ((~g4500));
assign g11024 = (g435&g10974);
assign g7058 = ((~II11255));
assign g11547 = ((~g11519));
assign g5904 = ((~II9539));
assign II14570 = ((~g9028));
assign II15368 = ((~g9990));
assign g7689 = ((~II12322));
assign II13908 = ((~g8526))|((~II13907));
assign II14549 = ((~g9262));
assign g5522 = (g1633&g4289);
assign g4190 = ((~II7387));
assign II12936 = ((~g7983));
assign g5897 = (g2204&g5354);
assign II17290 = ((~g11363))|((~II17288));
assign g11066 = ((~g10974));
assign g8346 = ((~II13418));
assign g6244 = (g2255&g5151);
assign II9491 = ((~g5072));
assign g7279 = ((~g6382));
assign II5218 = ((~g1104));
assign g8799 = (g8647&g8727);
assign II6145 = ((~g646))|((~II6143));
assign g10436 = ((~g10354)&(~g3566));
assign g7323 = ((~II11617));
assign g7318 = ((~II11602));
assign II16577 = ((~g10825));
assign g6453 = ((~g5817));
assign g8847 = ((~g8760))|((~g8683));
assign g5781 = (g1537&g5222);
assign II11656 = ((~g7122));
assign II17327 = ((~g11349));
assign II14418 = ((~g8941));
assign g11482 = (g6628)|(g11459);
assign II17173 = ((~g11293));
assign II12360 = ((~g7183));
assign gbuf14 = (g1356);
assign II7671 = ((~g3351));
assign II17710 = ((~g11620));
assign g10083 = ((~II15311));
assign g6786 = (g178&g5919);
assign g7980 = ((~II12786));
assign g8993 = ((~II14400));
assign g9745 = ((~g9454));
assign g4776 = ((~g3586));
assign g2435 = ((~g201));
assign g7819 = (g1887&g7479);
assign II11191 = ((~g6514));
assign g9412 = (g1727&g9052);
assign g7124 = ((~II11363));
assign g6928 = (g6359)|(g5703);
assign II16074 = ((~g10373))|((~II16072));
assign II7140 = ((~g2641));
assign g8632 = ((~II13915));
assign II11560 = ((~g7037));
assign g11166 = (g542&g11112);
assign II17359 = ((~g11372));
assign II11641 = ((~g6960));
assign g11458 = (g11426&g5446);
assign II13630 = ((~g8334));
assign II6611 = ((~g2626));
assign II15792 = ((~g10279));
assign g7704 = (g682&g7197);
assign g8715 = (g8416)|(g8687);
assign g8286 = (g8107)|(g7823);
assign g5190 = (g1245&g4716);
assign g11398 = ((~II17237));
assign g3731 = ((~II6911));
assign II14799 = ((~g9661));
assign II6876 = ((~g2956));
assign II10509 = ((~g786))|((~II10507));
assign g2501 = (g448)|(g452)|(g421)|(II5576);
assign g10486 = ((~II16095));
assign g8259 = (g8028)|(g7719);
assign g6835 = ((~II10885));
assign g7789 = ((~II12532));
assign II15305 = ((~g10001));
assign II8503 = ((~g4445));
assign g2871 = ((~II6013));
assign g9350 = ((~II14555));
assign g8292 = ((~II13230));
assign g9609 = (g907&g9205);
assign g6717 = ((~II10706));
assign g9428 = (g1756&g9030);
assign g11460 = (g11428&g5446);
assign g3121 = ((~g2462));
assign g4102 = ((~II7244));
assign II13002 = ((~g8045));
assign g10074 = ((~II15299));
assign g6047 = (g2017&g4977);
assign II5592 = ((~g1696))|((~II5591));
assign II15892 = ((~g10286))|((~II15890));
assign II15899 = ((~g857))|((~II15898));
assign II8919 = ((~g4576));
assign g8080 = ((~II12942));
assign II4850 = ((~g1958));
assign g5646 = ((~II9099));
assign g3987 = (g243&g3164);
assign g9855 = (g302&g9772);
assign g9082 = ((~g8892));
assign g11011 = (g1968&g10809);
assign g2764 = ((~II5850));
assign II16528 = ((~g10732));
assign II11456 = ((~g6440));
assign II5128 = ((~g1389))|((~II5126));
assign g4676 = ((~g3354));
assign g8078 = ((~II12936));
assign g4369 = ((~II7668));
assign g5124 = ((~g4596));
assign g10819 = ((~II16525));
assign II7468 = ((~g3697));
assign g8887 = (g8842)|(g8755);
assign II8298 = ((~g4437));
assign g5901 = ((~g5361));
assign g2528 = (g861)|(g857)|(g853)|(g849);
assign II12857 = ((~g7638));
assign II6565 = ((~g2614));
assign II8729 = ((~g4605))|((~II8728));
assign g7888 = (g7465&g7025);
assign g3427 = ((~g3144));
assign g8353 = ((~II13439));
assign g8217 = (g1872&g7883);
assign II13956 = ((~g8451));
assign g6944 = ((~II11082));
assign II14364 = ((~g8952));
assign g6290 = ((~II10129));
assign g9769 = ((~II14918));
assign II4903 = ((~g259));
assign g3765 = ((~g3120));
assign g8073 = (g709&g7826);
assign g8973 = (g8821)|(g8735);
assign g3070 = ((~g2016))|((~g1206));
assign g4523 = ((~g3546));
assign g10883 = ((~g10809));
assign g11226 = (g461&g11057);
assign g10344 = ((~II15798));
assign g5556 = ((~g4787)&(~g2695)&(~g2299)&(~g2031));
assign II8779 = ((~g4630))|((~II8778));
assign II8004 = ((~g3967));
assign II13574 = ((~g8360));
assign g11187 = (g5597&g11061);
assign g4384 = ((~II7707));
assign g8992 = ((~II14397));
assign g10196 = ((~II15562));
assign II16793 = ((~g11014));
assign II15406 = ((~g10065));
assign II9332 = ((~g4935));
assign II6370 = ((~g2356));
assign g7623 = (g664&g7079);
assign g11312 = (g11222)|(g11101);
assign g4320 = ((~g4013));
assign II6294 = ((~g2238));
assign g10171 = ((~II15507));
assign g7893 = (g7478&g7031);
assign g11427 = ((~II17334));
assign g7979 = ((~II12783));
assign g6585 = ((~II10541));
assign g4902 = (g1848&g4243);
assign g5175 = ((~g4682));
assign g9937 = (g9916&g9624);
assign II5116 = ((~g40));
assign g3009 = ((~g2135));
assign g7057 = ((~II11252));
assign g11497 = ((~II17510));
assign g6098 = (g1065&g5320);
assign g2840 = ((~II5960));
assign g10781 = ((~II16475));
assign II16148 = (g10386)|(g10384)|(g10476)|(g10474);
assign g9666 = ((~II14793));
assign g4281 = ((~g3586));
assign II6461 = ((~g2261));
assign II10299 = ((~g6243));
assign g5685 = ((~II9208));
assign g4360 = (g1861&g3748);
assign II15733 = ((~g10257));
assign g6538 = (g5782)|(g5006);
assign II8528 = ((~g4879))|((~II8527));
assign g4055 = ((~g3144));
assign II14101 = ((~g8774));
assign II15272 = ((~g10019));
assign II9759 = ((~g5344));
assign g10132 = ((~g10063));
assign g4754 = ((~g3440));
assign II11354 = ((~g6553));
assign g5557 = ((~g4538))|((~g3071))|((~g3011));
assign II10991 = ((~g6759));
assign g3088 = ((~II6294));
assign g3818 = ((~g3056))|((~g3071))|((~g2310))|((~g3003));
assign II11255 = ((~g6547));
assign g8230 = (g7515)|(g7991);
assign g10358 = ((~g10226)&(~g4620));
assign II10917 = ((~g6732));
assign g8221 = (g7496)|(g7993);
assign II16583 = ((~g10848));
assign g10476 = ((~II16038))|((~II16039));
assign g9880 = ((~g9751)&(~g9536)&(~g9557)&(~II15051));
assign g6027 = ((~g4566))|((~g4921));
assign g10444 = ((~g10325));
assign g9655 = ((~g9010)&(~g9240)&(~g9223)&(~II14776));
assign g7945 = (g2847&g7473);
assign II13538 = ((~g658))|((~II13537));
assign g10804 = ((~II16514));
assign g2942 = ((~II6121));
assign g3524 = ((~g3209))|((~g3221));
assign g2949 = ((~II6150));
assign g6526 = (g76&g6052);
assign g10909 = ((~II16679));
assign g2838 = ((~g2165));
assign g6548 = ((~g6132))|((~g6124))|((~g6122));
assign g6042 = (g5535)|(g3987);
assign g4554 = (g542&g3996);
assign g9759 = ((~g9454)&(~g9274)&(~g9292));
assign II5804 = (g2111)|(g2109)|(g2106)|(g2104);
assign g9530 = ((~II14675));
assign g11376 = (g11318&g4277);
assign g10371 = ((~g10344)&(~g3463));
assign II14607 = (g8995)|(g9205)|(g9192);
assign g6218 = ((~II9965));
assign g6916 = (g6348)|(g5687);
assign g4729 = ((~g3586));
assign II11309 = ((~g6531));
assign g6234 = (g2244&g5151);
assign g8440 = ((~II13618));
assign II9789 = ((~g5401));
assign II8479 = ((~g4455))|((~g3530));
assign g5013 = ((~g4749))|((~g3247))|((~g3205));
assign II6109 = ((~g2205))|((~g1494));
assign g8683 = (g4803&g8549);
assign g4544 = ((~g3880));
assign g4416 = ((~g3638));
assign g6791 = (g269&g5880);
assign g4576 = (g530&g4049);
assign II11752 = ((~g7032));
assign II16664 = ((~g10795));
assign g10623 = (g10544&g4536);
assign g9730 = (g9414)|(g9425)|(g9423);
assign g6180 = (g2190&g5128);
assign g7739 = (g6957&g3880);
assign II9766 = ((~g5348));
assign g5692 = ((~II9221));
assign g10465 = ((~II15986));
assign g4968 = (g1432&g4682);
assign g9268 = (g6681&g8947);
assign g11449 = ((~II17401))|((~II17402));
assign II5184 = ((~g1415))|((~g1515));
assign II11140 = ((~g6448));
assign g3292 = ((~g2373));
assign g8554 = (g8407&g8020);
assign g7378 = (g6990&g3880);
assign g8545 = ((~g3710))|((~g8390));
assign g2521 = (g538)|(g542)|(g476)|(II5626);
assign g8098 = (g6201&g7852);
assign g4390 = ((~g3914));
assign g2309 = (II5357)|(II5358);
assign g11243 = ((~g11112));
assign g5543 = (g4874&g4312);
assign II12805 = ((~g7684));
assign g7343 = ((~II11677));
assign g6478 = (g5706)|(g4967);
assign g7934 = ((~g7395))|((~g6847))|((~g7279))|((~g7369));
assign II15421 = ((~g10083));
assign II12843 = ((~g7683));
assign g10461 = ((~II15974));
assign g5255 = (g682&g4754);
assign II15341 = ((~g10019));
assign g8734 = (g8626&g7923);
assign g11301 = ((~II17084));
assign g5755 = (g5103&g5354);
assign II13308 = ((~g8190))|((~II13307));
assign II13809 = ((~g8480));
assign g11147 = (g321&g10929);
assign II17716 = ((~g11622));
assign g7917 = ((~g7497));
assign g10118 = ((~II15362));
assign II10840 = ((~g6719));
assign g11275 = (g11248)|(g11148);
assign g2109 = ((~II4996))|((~II4997));
assign g5266 = (g718&g4766);
assign II7916 = ((~g3664));
assign g6399 = ((~II10305));
assign II10114 = ((~g5768));
assign II14582 = (g8995)|(g9205)|(g9192);
assign II5754 = ((~g2304));
assign II6432 = ((~g2350));
assign g11252 = (g11099)|(g10969);
assign II11472 = ((~g6488));
assign II14944 = ((~g9454));
assign II9475 = ((~g5445));
assign g5229 = (g4364)|(g3516);
assign II11605 = ((~g6834));
assign II10663 = ((~g6040));
assign II7586 = ((~g4127));
assign II4869 = ((~g253));
assign II17424 = ((~g11424));
assign g6564 = ((~g5784));
assign g6403 = ((~g6128));
assign g4942 = ((~II8308));
assign g3461 = ((~II6671));
assign II13741 = ((~g8296));
assign g5007 = ((~II8379));
assign g6860 = ((~g6475));
assign II15350 = ((~g10001));
assign II15371 = ((~g9990));
assign g8773 = (g5491)|(g8653);
assign g7369 = ((~g7273));
assign II13825 = ((~g8488));
assign g10178 = ((~II15526));
assign g5023 = (g1071&g4511);
assign g2102 = ((~II4955))|((~II4956));
assign II5229 = ((~g182))|((~g148));
assign g5272 = ((~II8724));
assign g2478 = ((~g1610)&(~g1737));
assign II14188 = ((~g8792));
assign g11465 = (g11434&g5446);
assign g8326 = ((~II13360));
assign g4098 = ((~II7240));
assign g5144 = ((~g4682));
assign g6002 = (g5489)|(g3939);
assign g4615 = ((~II8024));
assign g7088 = (g2331&g6737);
assign g2937 = ((~II6106));
assign g6627 = (g58&g6181);
assign II7685 = ((~g3460))|((~II7683));
assign II9359 = ((~g5576));
assign II6760 = ((~g2943))|((~g1448));
assign II12271 = ((~g7218));
assign II17534 = ((~g11495));
assign g3061 = ((~g611))|((~g2374));
assign g5195 = ((~g4453));
assign II6844 = ((~g2915));
assign II14503 = ((~g8920));
assign g9505 = ((~g9052));
assign g3348 = ((~g2733));
assign II11716 = ((~g7026));
assign II9074 = ((~g4764));
assign g5063 = ((~g4363));
assign g6887 = (g6187&g6566);
assign II12942 = ((~g7982));
assign g8405 = ((~II13514))|((~II13515));
assign g7415 = ((~II11797));
assign g5998 = ((~II9620));
assign II8442 = ((~g4464));
assign g8950 = ((~II14303));
assign II13907 = ((~g8526))|((~g1432));
assign g2380 = ((~II5460))|((~II5461));
assign g7970 = (g7384&g7703);
assign g10595 = (g10550&g4347);
assign II8421 = ((~g4309));
assign g10388 = ((~g10305));
assign g7740 = (g7209)|(g6741);
assign g6948 = ((~II11088));
assign g5728 = ((~II9276));
assign g5320 = ((~g4418));
assign g6285 = ((~II10114));
assign g6638 = (g64&g6195);
assign g6811 = ((~II10843));
assign II10937 = ((~g6552));
assign g3069 = ((~II6277));
assign II13418 = ((~g8145));
assign g7116 = ((~II11351));
assign II12553 = ((~g7676));
assign II16292 = ((~g10551));
assign g11451 = ((~II17410));
assign g4836 = (g643&g3520);
assign g2348 = ((~II5418));
assign g8770 = (g5476)|(g8651);
assign II11997 = ((~g127))|((~II11995));
assign II17613 = ((~g11550));
assign g6192 = ((~II9923));
assign g6195 = ((~g5426));
assign II10825 = ((~g6588));
assign II14409 = ((~g8938));
assign g2080 = ((~II4894));
assign II9744 = ((~g5263));
assign g4586 = ((~g4089));
assign g7910 = ((~g7460));
assign g3714 = (g1690&g2991);
assign g5348 = ((~II8815));
assign g3411 = ((~II6616));
assign II17666 = ((~g11603));
assign g11317 = ((~II17112));
assign II13427 = ((~g8241));
assign g8726 = (g8608&g7913);
assign g6501 = (g5726)|(g4987);
assign g8093 = ((~II12948));
assign II7782 = ((~g3775));
assign II11498 = ((~g6578));
assign g8300 = ((~II13259))|((~II13260));
assign II5230 = ((~g182))|((~II5229));
assign g10184 = ((~g10039));
assign II9594 = ((~g5083));
assign g3439 = ((~g3144));
assign g3418 = (g2379&g3012);
assign g5493 = (g1923&g4265);
assign g5699 = (g1592&g5117);
assign g4344 = ((~g3946));
assign g7077 = ((~II11306));
assign g2224 = ((~g695));
assign II5949 = ((~g2540));
assign II13466 = ((~g8160));
assign g2341 = ((~II5403));
assign g11341 = ((~II17146));
assign g4330 = (g1163&g3693);
assign II12335 = ((~g7133));
assign g7580 = ((~II12056));
assign g9878 = ((~g9754)&(~g9536)&(~g9560)&(~II15045));
assign II5406 = ((~g898));
assign g10313 = ((~II15741));
assign g9949 = (g9929&g9392);
assign II6929 = ((~g2846));
assign g11283 = (g4966&g11205);
assign II17116 = ((~g11229));
assign g5534 = ((~g4545));
assign II17315 = ((~g11393));
assign g8337 = ((~II13391));
assign II14319 = ((~g8816));
assign g9423 = ((~g9052)&(~g9030));
assign g11417 = ((~II17302));
assign g8270 = (g7894)|(g3434);
assign g7333 = ((~II11647));
assign g10509 = ((~g10436))|((~g6023));
assign g3546 = ((~g3307));
assign g11294 = (g6576)|(g11210);
assign g8792 = ((~II14105));
assign g10767 = (g5500)|(g10681);
assign g7674 = (g7004&g3880);
assign g6161 = ((~II9886));
assign g10266 = ((~g10129));
assign g2912 = ((~II6085));
assign g10796 = ((~II16500));
assign II17707 = ((~g11619));
assign II4992 = ((~g1170));
assign g6061 = (g5204)|(g4);
assign g4773 = ((~II8133));
assign g10249 = ((~g10135));
assign II17274 = ((~g11389));
assign II10314 = ((~g6251));
assign g4976 = ((~g2310))|((~g4604))|((~g3807));
assign g9923 = (g9865)|(g9707);
assign g9510 = (g9125)|(g9111);
assign g5885 = ((~g5361));
assign II16030 = ((~g829))|((~g10368));
assign g10848 = ((~II16546));
assign II16206 = ((~g10453));
assign II6484 = ((~g2073));
assign II13023 = ((~g8050));
assign g11636 = (g11624&g7936);
assign II16009 = ((~g2689))|((~II16007));
assign II16673 = ((~g10782));
assign g6037 = ((~g3305)&(~g5614));
assign g4077 = ((~II7202));
assign g7300 = (g7139)|(g6326);
assign g2648 = ((~II5765));
assign g10257 = ((~g10197));
assign II13893 = ((~g8529))|((~g1436));
assign II14218 = ((~g605))|((~II14216));
assign g6852 = ((~II10914));
assign g5113 = ((~II8503));
assign II6071 = ((~g2269));
assign g8028 = (g7375&g7436);
assign g4462 = ((~II7825));
assign g3738 = ((~g3062));
assign II10362 = ((~g6224));
assign II10427 = ((~g5839));
assign II5060 = ((~g1191));
assign g11106 = ((~g10974));
assign II13274 = ((~g8158))|((~II13272));
assign g5097 = (g1786&g4603);
assign g3637 = ((~II6818));
assign g9699 = (g284&g9432);
assign II13424 = ((~g8200));
assign g6578 = ((~II10526));
assign g3908 = (g186&g3164);
assign II9706 = ((~g5221));
assign g8153 = (g7888)|(g6875);
assign g6918 = (g6358)|(g4252);
assign II15494 = ((~g10117));
assign g4442 = ((~g3638));
assign II11483 = ((~g6567));
assign g4084 = ((~g3119));
assign g3749 = ((~II6938));
assign g8411 = ((~II13538))|((~II13539));
assign II4965 = ((~g406))|((~II4964));
assign g2159 = ((~II5080));
assign g2449 = ((~g790));
assign II17362 = ((~g11376));
assign II15741 = ((~g10260));
assign II13782 = ((~g8515));
assign g5625 = (g1053&g4399);
assign II8050 = ((~g4089));
assign II17219 = ((~g11292));
assign II17767 = ((~g11648));
assign g8199 = (g7902)|(g7444);
assign g9024 = ((~II14409));
assign II15068 = ((~g9710));
assign II10296 = ((~g6242));
assign g3430 = ((~II6643));
assign g6935 = ((~II11065));
assign g8538 = ((~II13747));
assign g6633 = (g354&g6191);
assign g8805 = ((~II14136));
assign g7133 = (g6616)|(g3067);
assign g11648 = ((~II17746));
assign g2888 = ((~II6046));
assign II14567 = ((~g9027));
assign II12493 = ((~g7650));
assign II12448 = ((~g7530));
assign g11177 = (g511&g11112);
assign g5083 = (g3709&g4586);
assign g2247 = ((~II5258));
assign g11064 = ((~g10974));
assign g7478 = (g6884)|(g6423);
assign II14323 = ((~g8817));
assign g2317 = ((~g622));
assign II13606 = ((~g8311));
assign g6889 = (g1941&g6427);
assign II13819 = ((~g8488));
assign II11391 = ((~g6387));
assign II14191 = ((~g8795));
assign g9324 = (g8879&g5708);
assign II11680 = ((~g7064));
assign g10567 = (g10514)|(g7378);
assign II16778 = ((~g10891));
assign g2250 = ((~II5264))|((~II5265));
assign II7202 = ((~g2647));
assign g10116 = ((~II15356));
assign II6150 = ((~g2122));
assign II16850 = ((~g10905));
assign II14477 = ((~g8943));
assign g7515 = (g7148&g2855);
assign g8567 = ((~II13794));
assign II15562 = ((~g10098));
assign g4392 = (g3273&g3829);
assign II10762 = ((~g6127));
assign g10093 = ((~II15326));
assign II16025 = ((~g2701))|((~II16023));
assign g5911 = (g3322&g4977);
assign II8641 = ((~g4278))|((~II8640));
assign II8061 = ((~g3381));
assign g4089 = (g1959)|(g3318);
assign g9885 = (g9739)|(g9598)|(g9662)|(g9746);
assign II12523 = ((~g7421));
assign g7912 = ((~g7651));
assign II16283 = ((~g10538));
assign g10590 = ((~II16255));
assign g11303 = (g11214)|(g11092);
assign II11046 = ((~g6635));
assign g4473 = (g1125&g3874);
assign g5404 = (g4487)|(g3696);
assign g9535 = ((~II14690));
assign II5186 = ((~g1515))|((~II5184));
assign II12208 = ((~g7124));
assign g2040 = ((~g1786));
assign g3879 = ((~g3141)&(~g2354)&(~g2353));
assign II7694 = ((~g3742));
assign g2191 = ((~g1696));
assign II15210 = (g9839)|(g9964)|(g9852)|(g9882);
assign II14939 = ((~g9454));
assign II15114 = ((~g9875));
assign II15993 = ((~g10422))|((~II15992));
assign II16685 = ((~g10785));
assign g8751 = ((~g8632));
assign g5036 = (g4871)|(g4162);
assign g5647 = ((~II9102));
assign g8285 = (g8104)|(g7822);
assign g6891 = (g1950&g6435);
assign II10378 = ((~g6244));
assign II7043 = ((~g2908));
assign g10163 = ((~II15485));
assign g5501 = (g1672&g4273);
assign II10837 = ((~g6717));
assign g6808 = ((~II10834));
assign g3372 = ((~g3121));
assign g2481 = ((~g882));
assign g4176 = ((~II7345));
assign II13057 = ((~g7843));
assign g5844 = ((~II9461));
assign II8770 = ((~g4619))|((~g1133));
assign g4268 = ((~II7523));
assign g11173 = (g491&g11112);
assign II9114 = ((~g5603));
assign g6856 = ((~II10924));
assign g4747 = ((~g3586));
assign g2218 = ((~g85));
assign II10204 = ((~g6031));
assign g8085 = ((~g7932));
assign II5137 = ((~g525))|((~II5135));
assign g6246 = (g178&g5361);
assign g3254 = ((~g2322));
assign g5472 = ((~II8885));
assign g7072 = ((~II11293));
assign g8007 = ((~II12843));
assign II12565 = ((~g7388));
assign g10381 = ((~g10310)&(~g2998));
assign g8351 = ((~II13433));
assign g4890 = (g630&g4739);
assign g11044 = ((~II16793));
assign g9454 = (g8994&g5708);
assign g4581 = (g3766&g3254);
assign g3566 = ((~II6738));
assign g6418 = ((~g6137));
assign II12322 = ((~g7246));
assign g10891 = ((~II16635));
assign g6096 = (g5268)|(g4542);
assign g6831 = (g207&g6596);
assign g2863 = ((~g2316)&(~g2309));
assign g10198 = ((~II15568));
assign g4317 = ((~II7586));
assign II9084 = ((~g4886));
assign II14358 = ((~g8950));
assign g11082 = ((~II16859));
assign g8422 = ((~II13580));
assign II12040 = ((~g1466))|((~II12038));
assign g11429 = ((~II17340));
assign II8179 = ((~g3685))|((~II8178));
assign II12202 = ((~g6983));
assign g11553 = (g2683&g11519);
assign II12631 = ((~g7705));
assign g8988 = ((~II14385));
assign g7735 = ((~II12384));
assign II15299 = ((~g9995));
assign g6595 = ((~II10563));
assign II10613 = ((~g6000));
assign II17456 = ((~g11453));
assign g10336 = (g10230)|(g9572);
assign II12418 = ((~g7568));
assign II9296 = ((~g4908));
assign II13633 = ((~g8346));
assign g5483 = (g1621&g4254);
assign g5167 = ((~g4682));
assign g4787 = ((~g3423));
assign g2991 = ((~II6233));
assign g4602 = ((~II8011));
assign g10773 = (g5540)|(g10685);
assign g7027 = ((~II11176));
assign g10532 = ((~g10473));
assign II17540 = ((~g11498));
assign g3974 = (g231&g3164);
assign II6289 = ((~g981))|((~II6287));
assign II7810 = ((~g3799));
assign g5361 = (g4316)|(g4093)|(g126);
assign II9608 = ((~g5127));
assign II7746 = ((~g3763));
assign g7952 = ((~g7427));
assign II10910 = ((~g6703));
assign II6694 = ((~g2749));
assign g9826 = ((~II14979));
assign g9204 = ((~g6019))|((~g8942));
assign II17092 = ((~g11217));
assign II13887 = ((~g8532))|((~II13886));
assign g2200 = ((~g92));
assign g9770 = ((~g9432));
assign g11420 = ((~II17315));
assign g7435 = (g7260&g6572);
assign g7793 = ((~II12544));
assign g2257 = ((~II5283))|((~II5284));
assign g2169 = ((~g42));
assign II5461 = ((~g1003))|((~II5459));
assign g10445 = (g10315&g2135);
assign g6649 = ((~II10610));
assign g6209 = ((~II9956));
assign g5898 = ((~g5361));
assign g10285 = ((~g10276)&(~g3566));
assign g8279 = ((~II13209));
assign II16124 = ((~g10396));
assign g6304 = ((~II10171));
assign II6601 = ((~g3186));
assign II13788 = ((~g8517));
assign g10859 = (g5512)|(g10742);
assign II4979 = ((~g411))|((~II4978));
assign g3050 = ((~II6260));
assign II11734 = ((~g7024));
assign II10006 = ((~g5633));
assign g7811 = ((~II12598));
assign g8192 = ((~II13117));
assign g11323 = ((~II17124));
assign II17390 = ((~g11430));
assign g6653 = (g70&g6213);
assign g7919 = ((~g7512));
assign II8515 = ((~g3513))|((~II8513));
assign g2337 = ((~II5395));
assign g9110 = (g8880&g4790);
assign g7464 = ((~II11858));
assign g9266 = (g8932&g3398);
assign g2023 = ((~g1357));
assign g5539 = (g1684&g4314);
assign g4234 = ((~g3292)&(~g3793)&(~g2586)&(~g3776));
assign II11079 = ((~g6649));
assign g7471 = (g6880)|(g6416);
assign II13451 = ((~g8152));
assign g7762 = ((~II12451));
assign g10931 = ((~g10827));
assign g4288 = ((~g4130));
assign g3709 = ((~II6870));
assign g5640 = (g1059&g4427);
assign II12421 = ((~g7634));
assign g10057 = ((~II15278));
assign II5517 = ((~g1260))|((~II5516));
assign g8942 = ((~g8823))|((~g4921));
assign g4469 = ((~II7840));
assign g6292 = ((~II10135));
assign g11074 = ((~g10901));
assign g11091 = (g833&g10950);
assign g5891 = ((~g5361));
assign II9268 = ((~g5305));
assign g7771 = ((~II12478));
assign g4358 = (g1209&g3747);
assign g5588 = (g1639&g4508);
assign g4496 = ((~II7889));
assign g8927 = (g7872&g8807);
assign g9592 = (g4&g9292);
assign g3108 = (II6330&II6331);
assign g9589 = ((~g9125)&(~g9173)&(~g9151));
assign II15718 = ((~g10229))|((~II15716));
assign g5809 = (g5611)|(g4865);
assign g9668 = ((~g9490));
assign g7525 = ((~II11921));
assign g5783 = ((~II9377));
assign II11363 = ((~g6595));
assign g7559 = ((~II12009));
assign g6873 = (g3263&g6557);
assign II15829 = ((~g10203));
assign g2707 = ((~g2041));
assign g7272 = ((~II11519));
assign II10078 = ((~g5729));
assign g8650 = ((~II13933));
assign g7503 = (g6887)|(g6430);
assign g4892 = (g632&g4739);
assign II4911 = ((~g386))|((~II4910));
assign g7620 = ((~II12208));
assign g8465 = ((~g8289));
assign g6146 = ((~II9863));
assign g10946 = (g5225&g10827);
assign g6772 = (g6228&g722);
assign II10289 = ((~g6003));
assign g2154 = ((~II5067));
assign g8811 = (g7935)|(g8722);
assign II16432 = ((~g10702));
assign g11549 = ((~II17585))|((~II17586));
assign g4869 = (g1083&g3638);
assign g3694 = ((~II6851));
assign g7446 = ((~g7148));
assign II7166 = ((~g2620));
assign g7550 = ((~g6974));
assign II11103 = ((~g6667));
assign g4165 = ((~g3164));
assign g10211 = ((~II15583));
assign II9346 = ((~g5281));
assign g9359 = (g1308&g9173);
assign g9733 = ((~II14876));
assign II15238 = ((~g9974));
assign g9693 = (g275&g9432);
assign II17746 = ((~g11643));
assign g5490 = ((~II8911));
assign II15675 = ((~g10133));
assign II10177 = ((~g6103));
assign g6882 = ((~II10974));
assign II7022 = ((~g2941));
assign g8548 = ((~g8390));
assign g10673 = (g10580&g9450);
assign II12433 = ((~g7657));
assign g3305 = ((~II6474));
assign g7659 = ((~II12274));
assign II15224 = (g8174)|(g9908)|(g9937)|(g9834);
assign g3798 = ((~g3228));
assign II6316 = (g2082&g2087&g2381&g2395);
assign g10237 = (g10145&g9100);
assign g5616 = ((~II9046));
assign g7843 = (g7599&g5919);
assign g4242 = ((~g3664));
assign II10105 = ((~g5736));
assign g9356 = ((~II14573));
assign g1974 = ((~g627));
assign g2725 = ((~g2018));
assign g6030 = ((~II9639));
assign g9416 = ((~g9052)&(~g9030));
assign g7852 = ((~g7479));
assign g3388 = ((~II6590));
assign II14701 = ((~g9291));
assign g4260 = ((~II7513));
assign g11653 = ((~II17761));
assign g5000 = (g1470&g4640);
assign g8624 = ((~g8486));
assign II9988 = ((~g5526));
assign g9291 = ((~g8892));
assign II10949 = ((~g6747));
assign g4822 = ((~g3706));
assign g8136 = (g7926&g7045);
assign II7322 = ((~g3047))|((~II7321));
assign II6587 = ((~g2620));
assign g4867 = ((~II8204));
assign g9085 = ((~g8892));
assign g10120 = ((~II15368));
assign g8268 = (g7962)|(g7613);
assign g8838 = (g8602&g8702);
assign g4908 = ((~g4396));
assign g8103 = ((~g7994));
assign g8933 = ((~II14271))|((~II14272));
assign II12067 = ((~g7116))|((~g139));
assign II16039 = ((~g2707))|((~II16037));
assign II6200 = ((~g2525))|((~II6199));
assign II11707 = ((~g7009));
assign g10139 = ((~II15415));
assign g5354 = (g2733&g4460);
assign II6302 = ((~g2243));
assign g6833 = (g186&g6596);
assign II5540 = ((~g1023))|((~II5538));
assign g8705 = ((~II13991))|((~II13992));
assign II16356 = ((~g10597));
assign g6349 = ((~II10258));
assign g2809 = ((~II5909));
assign g8746 = ((~g8617))|((~g6517))|((~g6509));
assign g8731 = (g8622&g7918);
assign g5301 = ((~g4373));
assign g7798 = ((~II12559));
assign II15665 = ((~g10193));
assign g5596 = ((~II9020));
assign g11228 = (g466&g11060);
assign II9421 = ((~g5063));
assign g4529 = (g448&g3980);
assign g3727 = ((~II6901));
assign II17237 = ((~g11394));
assign g6411 = ((~g6135));
assign g8696 = ((~g8656));
assign g10539 = ((~II16184));
assign II7546 = ((~g4105));
assign g2540 = ((~II5655));
assign g2077 = ((~g219));
assign g9954 = (g9946)|(g9940)|(g9781);
assign g3012 = ((~II6247));
assign g3624 = ((~II6767));
assign g6539 = ((~II10461));
assign II8872 = ((~g4529));
assign II8465 = ((~g4807));
assign g2851 = ((~II5979));
assign g9780 = ((~g9474));
assign g11164 = (g4889&g11112);
assign II7952 = ((~g3664));
assign g2508 = ((~g940));
assign g9346 = ((~II14543));
assign g3910 = ((~g3015));
assign g7292 = (g7055)|(g6318);
assign g4224 = (g1092&g3638);
assign g7572 = ((~II12039))|((~II12040));
assign g6813 = ((~II10849));
assign II14232 = ((~g8800));
assign g4143 = ((~II7291));
assign g2304 = ((~II5348));
assign II8231 = ((~g4170));
assign g3793 = ((~g2593));
assign g6905 = ((~II11011));
assign g3219 = ((~II6395));
assign g6671 = (g342&g6227);
assign g3800 = ((~g3292));
assign g2948 = ((~II6144))|((~II6145));
assign II8109 = ((~g3622));
assign g6344 = ((~II10251));
assign II5418 = ((~g907));
assign II14394 = ((~g8884));
assign g3101 = (II6309&II6310);
assign g8506 = ((~g3475))|((~g8366));
assign g9910 = (g9892&g9809);
assign II9153 = ((~g5027));
assign g4223 = (g1003&g3914);
assign g10130 = ((~II15392));
assign g11282 = (g4958&g11203);
assign II15317 = ((~g10025));
assign g3998 = (g2677&g2276);
assign g5188 = (g4504&g4496);
assign g4886 = ((~II8231));
assign g4674 = ((~II8050));
assign g11576 = ((~II17610));
assign g4124 = ((~II7269));
assign II9108 = ((~g5593));
assign II13615 = ((~g8333));
assign II11746 = ((~g6857));
assign g6331 = (g201&g5904);
assign II10819 = ((~g6706));
assign g6104 = ((~II9769));
assign g3975 = ((~g3121));
assign g10488 = ((~II16101));
assign II16525 = ((~g10719));
assign g10129 = ((~II15389));
assign II6746 = ((~g2938))|((~g1453));
assign II11183 = ((~g6507));
assign II11901 = ((~g6897));
assign II12015 = ((~g6924));
assign g10683 = ((~g10612));
assign II10248 = ((~g6125));
assign g4215 = ((~II7462));
assign II5555 = ((~g110));
assign g6328 = (g1260&g5949);
assign II5276 = ((~g1411));
assign g6053 = ((~II9684));
assign g10788 = (g8303&g10754);
assign g11495 = ((~II17500));
assign g6043 = ((~II9662));
assign g7299 = (g7138)|(g6325);
assign II15184 = ((~g9974));
assign g4278 = ((~g3800)&(~g2593)&(~g2586)&(~g3776));
assign g5665 = ((~II9156));
assign g4431 = (g2268&g3533);
assign g7693 = ((~II12326));
assign g10322 = ((~g9317)&(~g10272));
assign II10855 = ((~g6685));
assign II5879 = ((~g2120))|((~II5878));
assign g11560 = (g2765&g11519);
assign g9814 = ((~g9490));
assign II15442 = ((~g10035))|((~II15441));
assign g8956 = ((~II14319));
assign II15437 = ((~g10050));
assign g5181 = (g4520&g4510);
assign g5317 = ((~II8796))|((~II8797));
assign g3204 = ((~g2571))|((~g2061));
assign II5880 = ((~g2115))|((~II5878));
assign g10933 = (g10853&g3982);
assign II10171 = ((~g5992));
assign g8262 = (g7970)|(g7625);
assign g2162 = ((~II5089));
assign g6354 = ((~g5867));
assign g7542 = (g7148&g2885);
assign g6072 = ((~g4977));
assign II7182 = ((~g2645));
assign II14602 = (g8995)|(g9205)|(g9192);
assign II15832 = ((~g10206));
assign g6016 = ((~II9632));
assign II5475 = ((~g1289));
assign g9952 = (g9944)|(g9938)|(g9817);
assign II7029 = ((~g2946));
assign g7618 = ((~II12202));
assign g6532 = (g339&g6057);
assign g2829 = ((~II5943));
assign g10734 = ((~II16413));
assign II12981 = ((~g8041));
assign g6757 = (g2221&g5919);
assign g4049 = ((~g3144));
assign g4782 = ((~g4089));
assign g2297 = ((~g865));
assign g4171 = ((~II7330));
assign II9712 = ((~g5230));
assign g4273 = ((~g4013));
assign g11641 = (g11615&g7901);
assign g2951 = (g2411&g1681);
assign II11662 = ((~g7033));
assign g7597 = ((~II12133));
assign g8126 = ((~II12989));
assign g5707 = (g1595&g5122);
assign g4166 = ((~II7315));
assign II12035 = ((~g6930));
assign g5938 = ((~g2764)&(~g4988));
assign II8473 = ((~g4577));
assign II11569 = ((~g6821));
assign g7257 = (g6701)|(g4725);
assign g5088 = ((~II8456));
assign g9604 = (g1194&g9111);
assign g6270 = ((~II10069));
assign g7414 = ((~II11794));
assign g5103 = ((~II8480))|((~II8481));
assign g4485 = ((~g3546));
assign II5435 = ((~g18));
assign II15971 = ((~g10408));
assign g4438 = ((~II7790));
assign g10873 = ((~II16589));
assign g8408 = (g704&g8139);
assign g9648 = (g16&g9274);
assign g5296 = ((~g4444));
assign g2605 = ((~II5716));
assign g7122 = ((~II11357));
assign g4875 = (g995&g3914);
assign II5704 = ((~g2056));
assign II11692 = ((~g7048));
assign II15204 = (g8168)|(g9904)|(g9933)|(g9829);
assign g9942 = (g9922&g9367);
assign II14614 = ((~g611))|((~II14612));
assign g3111 = (II6337&II6338);
assign g9984 = ((~II15184));
assign II5324 = ((~g1336))|((~II5323));
assign g8870 = ((~II14182));
assign g2031 = ((~g1690));
assign g6388 = ((~II10286));
assign g8920 = (g8845)|(g8759);
assign g9657 = (g919&g9205);
assign II14299 = ((~g8810));
assign II15430 = ((~g10047))|((~g10044));
assign g6581 = ((~II10531));
assign g3227 = ((~II6406));
assign II5571 = (g396)|(g391)|(g386)|(g426);
assign g5702 = ((~II9243));
assign II6133 = ((~g2253));
assign g6719 = ((~II10710));
assign g4557 = ((~g3946));
assign g3381 = (g940&g2756);
assign g7245 = (g6696)|(g6102);
assign g6749 = ((~II10756));
assign II6679 = ((~g2902));
assign II9138 = ((~g5210));
assign g6079 = (g1053&g5320);
assign II16053 = ((~g10371))|((~II16051));
assign g4381 = ((~g3914));
assign g7533 = ((~II11936))|((~II11937));
assign II13284 = ((~g1927))|((~II13283));
assign g2620 = ((~g1998));
assign II5824 = ((~g2502));
assign g8515 = ((~II13714));
assign II10810 = ((~g6539));
assign II9995 = ((~g5536));
assign g6845 = ((~II10907));
assign II17585 = ((~g11354))|((~II17584));
assign II14713 = ((~g9052));
assign g4112 = ((~g2994));
assign g8481 = ((~g8324));
assign g11198 = (g4919&g11069);
assign II5695 = ((~g575));
assign g6119 = ((~II9810));
assign II15701 = ((~g10236));
assign g10701 = (g10620&g10619);
assign g3979 = (g237&g3164);
assign II7054 = ((~g3093));
assign II17555 = ((~g11503));
assign II7224 = ((~g2981))|((~II7223));
assign II13485 = ((~g8194));
assign g9620 = (g2653&g9240);
assign g8498 = ((~g8353));
assign g11025 = (g426&g10974);
assign g2638 = ((~II5751));
assign g2197 = ((~g101));
assign g7759 = ((~II12442));
assign g2756 = (g936&g2081);
assign g4680 = ((~g3829));
assign g4450 = ((~g3914));
assign II15075 = ((~g9761));
assign g10240 = (g10150&g9103);
assign II16037 = ((~g10427))|((~g2707));
assign II9773 = ((~g4934));
assign II9180 = ((~g4905));
assign g5942 = ((~II9575))|((~II9576));
assign g8947 = (g8056&g6368&g8828);
assign II5445 = ((~g922));
assign II13965 = ((~g8451));
assign g2779 = ((~g1974));
endmodule
